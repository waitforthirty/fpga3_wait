
#******
# Preview export LEF
#
#	 Preview sub-version 5.10.41.500.5.95
#
# REF LIBS: myvtvt_tsmc180_lib 
# TECH LIB NAME: dump_tsmc180_techlib
# TECH FILE NAME: techfile.cds
#******

VERSION 5.5 ;

NAMESCASESENSITIVE ON ;

DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

UNITS
    DATABASE MICRONS 1000  ;
END UNITS

 MANUFACTURINGGRID    0.045000 ;
LAYER nwell
    TYPE MASTERSLICE ;
END nwell

LAYER nactive
    TYPE MASTERSLICE ;
END nactive

LAYER pactive
    TYPE MASTERSLICE ;
END pactive

LAYER poly
    TYPE MASTERSLICE ;
END poly

LAYER glass
    TYPE MASTERSLICE ;
END glass

LAYER pad
    TYPE MASTERSLICE ;
END pad

LAYER sblock
    TYPE MASTERSLICE ;
END sblock

LAYER text
    TYPE MASTERSLICE ;
END text

LAYER res_id
    TYPE MASTERSLICE ;
END res_id

LAYER cap_id
    TYPE MASTERSLICE ;
END cap_id

LAYER metalcap
    TYPE MASTERSLICE ;
END metalcap

LAYER nodrc
    TYPE MASTERSLICE ;
END nodrc

LAYER cc
    TYPE CUT ;
    SPACING 0.360 ;
END cc

LAYER metal1
    TYPE ROUTING ;
    WIDTH 0.270 ;
    SPACING 0.270 ;
    OFFSET 0.000 ;
    PITCH 0.810 ;
    DIRECTION HORIZONTAL ;
    CAPACITANCE CPERSQDIST 38.0000000000 ;
    RESISTANCE RPERSQ 0.08000000 ;
END metal1

LAYER via
    TYPE CUT ;
    SPACING 0.270 ;
END via

LAYER metal2
    TYPE ROUTING ;
    WIDTH 0.270 ;
    SPACING 0.360 ;
    OFFSET 0.000 ;
    PITCH 0.810 ;
    DIRECTION VERTICAL ;
    CAPACITANCE CPERSQDIST 18.0000000000 ;
    RESISTANCE RPERSQ 0.08000000 ;
END metal2

LAYER via2
    TYPE CUT ;
    SPACING 0.270 ;
END via2

LAYER metal3
    TYPE ROUTING ;
    WIDTH 0.270 ;
    SPACING 0.360 ;
    OFFSET 0.000 ;
    PITCH 0.810 ;
    DIRECTION HORIZONTAL ;
    CAPACITANCE CPERSQDIST 13.0000000000 ;
    RESISTANCE RPERSQ 0.08000000 ;
END metal3

LAYER via3
    TYPE CUT ;
    SPACING 0.360 ;
END via3

LAYER metal4
    TYPE ROUTING ;
    WIDTH 0.270 ;
    SPACING 0.360 ;
    OFFSET 0.000 ;
    PITCH 0.810 ;
    DIRECTION VERTICAL ;
    CAPACITANCE CPERSQDIST 8.0000000000 ;
    RESISTANCE RPERSQ 0.08000000 ;
END metal4

LAYER via4
    TYPE CUT ;
    SPACING 0.270 ;
END via4

LAYER metal5
    TYPE ROUTING ;
    WIDTH 0.360 ;
    SPACING 0.360 ;
    OFFSET 0.000 ;
    PITCH 0.810 ;
    DIRECTION HORIZONTAL ;
    CAPACITANCE CPERSQDIST 8.0000000000 ;
    RESISTANCE RPERSQ 0.07000000 ;
END metal5

LAYER via5
    TYPE CUT ;
    SPACING 0.360 ;
END via5

LAYER metal6
    TYPE ROUTING ;
    WIDTH 0.450 ;
    SPACING 0.450 ;
    OFFSET 0.000 ;
    PITCH 1.620 ;
    DIRECTION VERTICAL ;
    CAPACITANCE CPERSQDIST 3.0000000000 ;
    RESISTANCE RPERSQ 0.03000000 ;
END metal6

VIA M1_P
    LAYER pactive ;
        RECT -0.180 -0.180 0.180 0.180 ;
    LAYER cc ;
        RECT -0.090 -0.090 0.090 0.090 ;
    LAYER metal1 ;
        RECT -0.180 -0.180 0.180 0.180 ;
END M1_P

VIA M1_N
    LAYER nactive ;
        RECT -0.180 -0.180 0.180 0.180 ;
    LAYER cc ;
        RECT -0.090 -0.090 0.090 0.090 ;
    LAYER metal1 ;
        RECT -0.180 -0.180 0.180 0.180 ;
END M1_N

VIA NTAP
    LAYER nwell ;
        RECT -0.450 -0.450 0.450 0.450 ;
    LAYER cc ;
        RECT -0.090 -0.090 0.090 0.090 ;
    LAYER metal1 ;
        RECT -0.180 -0.180 0.180 0.180 ;
END NTAP

VIA M1_POLY
    LAYER poly ;
        RECT -0.180 -0.180 0.180 0.180 ;
    LAYER cc ;
        RECT -0.090 -0.090 0.090 0.090 ;
    LAYER metal1 ;
        RECT -0.180 -0.180 0.180 0.180 ;
END M1_POLY

VIA M2_M1 DEFAULT
    LAYER metal1 ;
        RECT -0.225 -0.225 0.225 0.225 ;
    LAYER via ;
        RECT -0.135 -0.135 0.135 0.135 ;
    LAYER metal2 ;
        RECT -0.225 -0.225 0.225 0.225 ;
END M2_M1

VIA M6_M5 DEFAULT
    LAYER metal5 ;
        RECT -0.315 -0.315 0.315 0.315 ;
    LAYER via5 ;
        RECT -0.225 -0.225 0.225 0.225 ;
    LAYER metal6 ;
        RECT -0.405 -0.405 0.405 0.405 ;
END M6_M5

VIA M5_M4 DEFAULT
    LAYER metal4 ;
        RECT -0.225 -0.225 0.225 0.225 ;
    LAYER via4 ;
        RECT -0.135 -0.135 0.135 0.135 ;
    LAYER metal5 ;
        RECT -0.225 -0.225 0.225 0.225 ;
END M5_M4

VIA M4_M3 DEFAULT
    LAYER metal3 ;
        RECT -0.225 -0.225 0.225 0.225 ;
    LAYER via3 ;
        RECT -0.135 -0.135 0.135 0.135 ;
    LAYER metal4 ;
        RECT -0.225 -0.225 0.225 0.225 ;
END M4_M3

VIA M3_M2 DEFAULT
    LAYER metal2 ;
        RECT -0.225 -0.225 0.225 0.225 ;
    LAYER via2 ;
        RECT -0.135 -0.135 0.135 0.135 ;
    LAYER metal3 ;
        RECT -0.225 -0.225 0.225 0.225 ;
END M3_M2

VIARULE viagen21 GENERATE
    LAYER metal1 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.090 ;
        METALOVERHANG 0.000 ;

    LAYER metal2 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.090 ;
        METALOVERHANG 0.000 ;

    LAYER via ;
        RECT -0.135 -0.135 0.135 0.135 ;
        SPACING 0.720 BY 0.720 ;
END viagen21

VIARULE viagen65 GENERATE
    LAYER metal5 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.090 ;
        METALOVERHANG 0.000 ;

    LAYER metal6 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.090 ;
        METALOVERHANG 0.000 ;

    LAYER via5 ;
        RECT -0.135 -0.135 0.135 0.135 ;
        SPACING 1.080 BY 1.080 ;
END viagen65

VIARULE viagen54 GENERATE
    LAYER metal5 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.090 ;
        METALOVERHANG 0.000 ;

    LAYER metal4 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.090 ;
        METALOVERHANG 0.000 ;

    LAYER via4 ;
        RECT -0.135 -0.135 0.135 0.135 ;
        SPACING 0.720 BY 0.720 ;
END viagen54

VIARULE viagen43 GENERATE
    LAYER metal3 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.090 ;
        METALOVERHANG 0.000 ;

    LAYER metal4 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.090 ;
        METALOVERHANG 0.000 ;

    LAYER via3 ;
        RECT -0.135 -0.135 0.135 0.135 ;
        SPACING 0.720 BY 0.720 ;
END viagen43

VIARULE viagen32 GENERATE
    LAYER metal3 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.090 ;
        METALOVERHANG 0.000 ;

    LAYER metal2 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.090 ;
        METALOVERHANG 0.000 ;

    LAYER via2 ;
        RECT -0.135 -0.135 0.135 0.135 ;
        SPACING 0.720 BY 0.720 ;
END viagen32

SITE CoreSite
    SYMMETRY Y  ;
    CLASS CORE  ;
    SIZE 0.810 BY 11.340 ;
END CoreSite

MACRO xor2_2
    CLASS CORE ;
    FOREIGN xor2_2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.290 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.860 4.680 5.985 5.040 ;
        RECT  4.275 5.490 5.220 5.850 ;
        RECT  4.860 3.870 5.220 5.850 ;
        RECT  4.230 3.870 5.220 4.230 ;
        RECT  4.275 5.490 4.635 9.270 ;
        RECT  4.230 2.160 4.590 4.230 ;
        END
    END op
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  6.345 6.345 6.615 6.615 ;
        RECT  2.295 6.345 2.565 6.615 ;
        LAYER metal2 ;
        RECT  6.255 6.255 6.705 6.705 ;
        RECT  2.205 6.300 6.705 6.660 ;
        RECT  2.205 6.255 2.655 6.705 ;
        LAYER metal1 ;
        RECT  6.255 6.255 6.705 6.705 ;
        RECT  2.205 6.255 2.655 6.705 ;
        END
    END ip1
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  4.230 4.725 4.500 4.995 ;
        RECT  0.675 4.725 0.945 4.995 ;
        LAYER metal2 ;
        RECT  4.140 4.635 4.590 5.085 ;
        RECT  0.585 4.680 4.590 5.040 ;
        RECT  0.585 4.635 1.035 5.085 ;
        LAYER metal1 ;
        RECT  4.140 4.635 4.590 5.085 ;
        RECT  0.585 4.635 1.035 5.085 ;
        END
    END ip2
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 7.290 11.340 ;
        RECT  5.535 6.750 5.895 11.340 ;
        RECT  2.970 7.785 3.330 11.340 ;
        RECT  0.630 6.750 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 7.290 0.990 ;
        RECT  5.535 0.000 5.895 3.420 ;
        RECT  2.970 0.000 3.330 3.420 ;
        RECT  0.630 0.000 0.990 3.420 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  1.395 5.445 1.845 5.895 ;
        RECT  1.440 2.160 1.800 9.270 ;
        RECT  3.015 3.825 3.465 4.275 ;
        RECT  3.060 3.825 3.420 5.040 ;
        RECT  2.250 4.680 3.420 5.040 ;
        RECT  2.250 2.160 2.610 5.850 ;
        RECT  2.250 5.490 3.420 5.850 ;
        RECT  3.060 5.490 3.420 7.425 ;
        RECT  2.250 7.065 3.420 7.425 ;
        RECT  2.250 7.065 2.610 9.270 ;
        RECT  5.580 5.445 6.030 5.895 ;
        RECT  6.255 3.825 6.705 4.275 ;
        LAYER via ;
        RECT  1.485 5.535 1.755 5.805 ;
        RECT  3.105 3.915 3.375 4.185 ;
        RECT  5.670 5.535 5.940 5.805 ;
        RECT  6.345 3.915 6.615 4.185 ;
        LAYER metal2 ;
        RECT  1.395 5.490 6.030 5.850 ;
        RECT  1.395 5.445 1.845 5.895 ;
        RECT  5.580 5.445 6.030 5.895 ;
        RECT  3.015 3.870 6.705 4.230 ;
        RECT  3.015 3.825 3.465 4.275 ;
        RECT  6.255 3.825 6.705 4.275 ;
    END
END xor2_2

MACRO xor2_1
    CLASS CORE ;
    FOREIGN xor2_1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.290 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  5.985 6.345 6.255 6.615 ;
        RECT  2.295 6.345 2.565 6.615 ;
        LAYER metal2 ;
        RECT  5.895 6.255 6.345 6.705 ;
        RECT  2.205 6.300 6.345 6.660 ;
        RECT  2.205 6.255 2.655 6.705 ;
        LAYER metal1 ;
        RECT  5.895 6.255 6.345 6.705 ;
        RECT  2.205 6.255 2.655 6.705 ;
        END
    END ip1
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  4.185 5.535 4.455 5.805 ;
        RECT  0.675 5.535 0.945 5.805 ;
        LAYER metal2 ;
        RECT  4.095 5.445 4.545 5.895 ;
        RECT  0.585 5.490 4.545 5.850 ;
        RECT  0.585 5.445 1.035 5.895 ;
        LAYER metal1 ;
        RECT  4.095 5.445 4.545 5.895 ;
        RECT  0.585 5.445 1.035 5.895 ;
        END
    END ip2
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.995 5.490 5.895 5.850 ;
        RECT  4.275 7.110 5.355 7.470 ;
        RECT  4.995 3.870 5.355 7.470 ;
        RECT  4.230 3.870 5.355 4.230 ;
        RECT  4.275 7.110 4.635 9.270 ;
        RECT  4.230 2.160 4.590 4.230 ;
        END
    END op
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 7.290 11.340 ;
        RECT  5.535 8.010 5.895 11.340 ;
        RECT  2.970 8.010 3.330 11.340 ;
        RECT  0.630 8.010 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 7.290 0.990 ;
        RECT  5.535 0.000 5.895 2.790 ;
        RECT  2.970 0.000 3.330 2.790 ;
        RECT  0.630 0.000 0.990 2.790 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  1.395 4.635 1.845 5.085 ;
        RECT  1.440 2.160 1.800 9.270 ;
        RECT  2.250 2.160 2.610 3.510 ;
        RECT  2.250 3.150 3.780 3.510 ;
        RECT  3.375 3.825 3.825 4.275 ;
        RECT  3.420 3.150 3.780 7.650 ;
        RECT  2.250 7.290 3.780 7.650 ;
        RECT  2.250 7.290 2.610 9.270 ;
        RECT  5.805 4.635 6.255 5.085 ;
        RECT  5.895 3.825 6.345 4.275 ;
        LAYER via ;
        RECT  1.485 4.725 1.755 4.995 ;
        RECT  3.465 3.915 3.735 4.185 ;
        RECT  5.895 4.725 6.165 4.995 ;
        RECT  5.985 3.915 6.255 4.185 ;
        LAYER metal2 ;
        RECT  1.395 4.680 6.255 5.040 ;
        RECT  1.395 4.635 1.845 5.085 ;
        RECT  5.805 4.635 6.255 5.085 ;
        RECT  3.375 3.870 6.345 4.230 ;
        RECT  3.375 3.825 3.825 4.275 ;
        RECT  5.895 3.825 6.345 4.275 ;
    END
END xor2_1

MACRO xnor2_2
    CLASS CORE ;
    FOREIGN xnor2_2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.100 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  5.715 6.345 5.985 6.615 ;
        RECT  2.295 6.345 2.565 6.615 ;
        LAYER metal2 ;
        RECT  5.625 6.255 6.075 6.705 ;
        RECT  2.205 6.300 6.075 6.660 ;
        RECT  2.205 6.255 2.655 6.705 ;
        LAYER metal1 ;
        RECT  5.625 6.255 6.075 6.705 ;
        RECT  2.205 6.255 2.655 6.705 ;
        END
    END ip1
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  4.140 4.725 4.410 4.995 ;
        RECT  0.675 4.725 0.945 4.995 ;
        LAYER metal2 ;
        RECT  4.050 4.635 4.500 5.085 ;
        RECT  0.585 4.680 4.500 5.040 ;
        RECT  0.585 4.635 1.035 5.085 ;
        LAYER metal1 ;
        RECT  4.050 4.635 4.500 5.085 ;
        RECT  0.585 4.635 1.035 5.085 ;
        END
    END ip2
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.110 6.300 7.470 9.270 ;
        RECT  6.615 3.870 7.470 4.230 ;
        RECT  7.110 2.160 7.470 4.230 ;
        RECT  6.615 6.300 7.470 6.660 ;
        RECT  6.615 3.870 6.975 6.660 ;
        END
    END op
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 8.100 11.340 ;
        RECT  6.300 6.975 6.660 11.340 ;
        RECT  5.490 8.010 5.850 11.340 ;
        RECT  2.880 8.010 3.240 11.340 ;
        RECT  0.630 8.010 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 8.100 0.990 ;
        RECT  6.300 0.000 6.660 3.420 ;
        RECT  5.490 0.000 5.850 2.790 ;
        RECT  2.880 0.000 3.240 2.790 ;
        RECT  0.630 0.000 0.990 2.790 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  1.395 5.445 1.845 5.895 ;
        RECT  1.440 2.160 1.800 9.270 ;
        RECT  2.160 2.160 2.520 3.420 ;
        RECT  2.160 3.060 3.735 3.420 ;
        RECT  3.330 3.825 3.780 4.275 ;
        RECT  3.375 3.060 3.735 7.470 ;
        RECT  2.160 7.110 3.735 7.470 ;
        RECT  2.160 7.110 2.520 9.270 ;
        RECT  5.625 3.825 6.075 4.275 ;
        RECT  4.140 2.160 4.500 3.420 ;
        RECT  4.140 3.060 5.355 3.420 ;
        RECT  4.995 4.680 6.165 5.040 ;
        RECT  4.995 3.060 5.355 6.210 ;
        RECT  4.185 5.850 5.355 6.210 ;
        RECT  4.185 5.850 4.545 9.270 ;
        RECT  5.805 5.445 6.255 5.895 ;
        LAYER via ;
        RECT  1.485 5.535 1.755 5.805 ;
        RECT  3.420 3.915 3.690 4.185 ;
        RECT  5.715 3.915 5.985 4.185 ;
        RECT  5.895 5.535 6.165 5.805 ;
        LAYER metal2 ;
        RECT  3.330 3.870 6.075 4.230 ;
        RECT  3.330 3.825 3.780 4.275 ;
        RECT  5.625 3.825 6.075 4.275 ;
        RECT  1.350 5.490 6.255 5.850 ;
        RECT  1.395 5.445 1.845 5.895 ;
        RECT  5.805 5.445 6.255 5.895 ;
    END
END xnor2_2

MACRO xnor2_1
    CLASS CORE ;
    FOREIGN xnor2_1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.100 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  5.715 6.345 5.985 6.615 ;
        RECT  2.295 6.345 2.565 6.615 ;
        LAYER metal2 ;
        RECT  5.625 6.255 6.075 6.705 ;
        RECT  2.205 6.300 6.075 6.660 ;
        RECT  2.205 6.255 2.655 6.705 ;
        LAYER metal1 ;
        RECT  5.625 6.255 6.075 6.705 ;
        RECT  2.205 6.255 2.655 6.705 ;
        END
    END ip1
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  4.140 4.725 4.410 4.995 ;
        RECT  0.675 4.725 0.945 4.995 ;
        LAYER metal2 ;
        RECT  4.050 4.635 4.500 5.085 ;
        RECT  0.585 4.680 4.500 5.040 ;
        RECT  0.585 4.635 1.035 5.085 ;
        LAYER metal1 ;
        RECT  4.050 4.635 4.500 5.085 ;
        RECT  0.585 4.635 1.035 5.085 ;
        END
    END ip2
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.110 6.300 7.470 9.270 ;
        RECT  6.615 3.870 7.470 4.230 ;
        RECT  7.110 2.160 7.470 4.230 ;
        RECT  6.615 6.300 7.470 6.660 ;
        RECT  6.615 3.870 6.975 6.660 ;
        END
    END op
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 8.100 11.340 ;
        RECT  6.300 8.010 6.660 11.340 ;
        RECT  5.490 8.010 5.850 11.340 ;
        RECT  2.880 8.010 3.240 11.340 ;
        RECT  0.630 8.010 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 8.100 0.990 ;
        RECT  6.300 0.000 6.660 2.790 ;
        RECT  5.490 0.000 5.850 2.790 ;
        RECT  2.880 0.000 3.240 2.790 ;
        RECT  0.630 0.000 0.990 2.790 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  1.395 5.445 1.845 5.895 ;
        RECT  1.440 2.160 1.800 9.270 ;
        RECT  2.160 2.160 2.520 3.420 ;
        RECT  2.160 3.060 3.735 3.420 ;
        RECT  3.330 3.825 3.780 4.275 ;
        RECT  3.375 3.060 3.735 7.470 ;
        RECT  2.160 7.110 3.735 7.470 ;
        RECT  2.160 7.110 2.520 9.270 ;
        RECT  5.625 3.825 6.075 4.275 ;
        RECT  4.140 2.160 4.500 3.420 ;
        RECT  4.140 3.060 5.355 3.420 ;
        RECT  4.995 4.680 6.165 5.040 ;
        RECT  4.995 3.060 5.355 6.210 ;
        RECT  4.185 5.850 5.355 6.210 ;
        RECT  4.185 5.850 4.545 9.270 ;
        RECT  5.805 5.445 6.255 5.895 ;
        LAYER via ;
        RECT  1.485 5.535 1.755 5.805 ;
        RECT  3.420 3.915 3.690 4.185 ;
        RECT  5.715 3.915 5.985 4.185 ;
        RECT  5.895 5.535 6.165 5.805 ;
        LAYER metal2 ;
        RECT  3.330 3.870 6.075 4.230 ;
        RECT  3.330 3.825 3.780 4.275 ;
        RECT  5.625 3.825 6.075 4.275 ;
        RECT  1.350 5.490 6.255 5.850 ;
        RECT  1.395 5.445 1.845 5.895 ;
        RECT  5.805 5.445 6.255 5.895 ;
    END
END xnor2_1

MACRO or4_4
    CLASS CORE ;
    FOREIGN or4_4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.480 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip4
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  3.870 5.445 4.230 5.805 ;
        END
    END ip4
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.860 3.870 5.220 6.480 ;
        RECT  4.680 2.160 5.040 4.230 ;
        RECT  4.545 6.120 4.905 9.270 ;
        END
    END op
    PIN ip3
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 4.680 2.610 5.040 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 5.490 1.800 5.850 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 6.300 0.990 6.660 ;
        END
    END ip1
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 6.480 11.340 ;
        RECT  5.310 6.750 5.670 11.340 ;
        RECT  3.825 6.750 4.185 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 6.480 0.990 ;
        RECT  5.400 0.000 5.760 3.420 ;
        RECT  3.870 0.000 4.230 3.420 ;
        RECT  2.250 0.000 2.610 3.420 ;
        RECT  0.630 0.000 0.990 3.420 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  1.440 2.160 1.800 4.230 ;
        RECT  1.440 3.870 3.420 4.230 ;
        RECT  3.060 4.500 4.410 4.860 ;
        RECT  3.060 2.160 3.420 6.660 ;
        RECT  1.485 6.300 3.420 6.660 ;
        RECT  1.485 6.300 1.845 9.270 ;
    END
END or4_4

MACRO or4_2
    CLASS CORE ;
    FOREIGN or4_2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.680 2.160 5.040 6.660 ;
        RECT  4.545 6.300 4.905 9.270 ;
        END
    END op
    PIN ip4
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  3.870 5.490 4.230 5.850 ;
        END
    END ip4
    PIN ip3
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 4.680 2.610 5.040 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 5.490 1.800 5.850 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 6.300 0.990 6.660 ;
        END
    END ip1
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 5.670 0.990 ;
        RECT  3.870 0.000 4.230 3.420 ;
        RECT  2.250 0.000 2.610 3.420 ;
        RECT  0.630 0.000 0.990 3.420 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 5.670 11.340 ;
        RECT  3.825 6.750 4.185 11.340 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  1.440 2.160 1.800 4.230 ;
        RECT  1.440 3.870 3.420 4.230 ;
        RECT  3.060 4.500 4.410 4.860 ;
        RECT  3.060 2.160 3.420 6.660 ;
        RECT  1.485 6.300 3.420 6.660 ;
        RECT  1.485 6.300 1.845 9.270 ;
    END
END or4_2

MACRO or4_1
    CLASS CORE ;
    FOREIGN or4_1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.680 2.160 5.040 7.470 ;
        RECT  4.545 7.110 4.905 9.270 ;
        END
    END op
    PIN ip4
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  3.060 4.680 3.420 5.040 ;
        END
    END ip4
    PIN ip3
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 5.490 2.610 5.850 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 6.300 1.800 6.660 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 3.060 0.990 3.420 ;
        END
    END ip1
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 5.670 0.990 ;
        RECT  3.870 0.000 4.230 2.790 ;
        RECT  2.250 0.000 2.610 2.790 ;
        RECT  0.630 0.000 0.990 2.790 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 5.670 11.340 ;
        RECT  3.825 8.010 4.185 11.340 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  2.205 6.255 2.655 6.705 ;
        RECT  2.250 6.255 2.610 7.470 ;
        RECT  1.485 7.110 2.610 7.470 ;
        RECT  1.485 7.110 1.845 9.270 ;
        RECT  1.440 2.160 1.800 3.420 ;
        RECT  1.440 3.060 3.420 3.420 ;
        RECT  3.060 2.160 3.420 4.230 ;
        RECT  3.060 3.870 4.230 4.230 ;
        RECT  3.870 3.870 4.230 6.705 ;
        RECT  3.825 6.255 4.275 6.705 ;
        LAYER via ;
        RECT  2.295 6.345 2.565 6.615 ;
        RECT  3.915 6.345 4.185 6.615 ;
        LAYER metal2 ;
        RECT  2.205 6.300 4.275 6.660 ;
        RECT  2.205 6.255 2.655 6.705 ;
        RECT  3.825 6.255 4.275 6.705 ;
    END
END or4_1

MACRO or3_4
    CLASS CORE ;
    FOREIGN or3_4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.480 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip3
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  3.060 3.870 3.420 4.230 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 4.680 2.610 5.040 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip1
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.005 2.160 4.365 3.780 ;
        RECT  3.465 4.680 4.230 5.040 ;
        RECT  3.870 3.420 4.230 5.040 ;
        RECT  3.465 4.680 3.825 9.270 ;
        END
    END op
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 6.480 11.340 ;
        RECT  4.275 6.750 4.635 11.340 ;
        RECT  2.610 6.750 2.970 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 6.480 0.990 ;
        RECT  4.815 0.000 5.175 3.420 ;
        RECT  3.195 0.000 3.555 3.420 ;
        RECT  1.575 0.000 1.935 3.150 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  0.765 2.160 1.125 3.780 ;
        RECT  2.385 2.160 2.745 3.780 ;
        RECT  0.765 3.420 2.745 3.780 ;
        RECT  1.530 5.445 1.980 5.895 ;
        RECT  1.575 3.420 1.935 6.660 ;
        RECT  0.765 6.300 1.935 6.660 ;
        RECT  0.765 6.300 1.125 9.270 ;
        RECT  4.590 5.445 5.040 5.895 ;
        LAYER via ;
        RECT  1.620 5.535 1.890 5.805 ;
        RECT  4.680 5.535 4.950 5.805 ;
        LAYER metal2 ;
        RECT  1.530 5.490 5.040 5.850 ;
        RECT  1.530 5.445 1.980 5.895 ;
        RECT  4.590 5.445 5.040 5.895 ;
    END
END or3_4

MACRO or3_2
    CLASS CORE ;
    FOREIGN or3_2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 4.680 1.800 5.040 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip1
    PIN ip3
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  3.060 3.870 3.420 4.230 ;
        END
    END ip3
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.005 2.160 4.365 3.780 ;
        RECT  2.835 4.680 4.230 5.040 ;
        RECT  3.870 3.420 4.230 5.040 ;
        RECT  3.465 6.165 3.825 9.270 ;
        RECT  2.835 6.165 3.825 6.525 ;
        RECT  2.835 4.680 3.195 6.525 ;
        END
    END op
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 5.670 0.990 ;
        RECT  3.195 0.000 3.555 3.420 ;
        RECT  1.575 0.000 1.935 3.150 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 5.670 11.340 ;
        RECT  2.610 6.795 2.970 11.340 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  0.765 2.160 1.125 3.780 ;
        RECT  2.385 2.160 2.745 3.780 ;
        RECT  0.765 3.420 2.745 3.780 ;
        RECT  2.070 3.420 2.430 5.895 ;
        RECT  1.980 5.445 2.430 5.895 ;
        RECT  1.665 5.490 2.025 6.750 ;
        RECT  0.765 6.390 2.025 6.750 ;
        RECT  0.765 6.390 1.125 9.270 ;
        RECT  3.510 5.445 3.960 5.895 ;
        LAYER via ;
        RECT  2.070 5.535 2.340 5.805 ;
        RECT  3.600 5.535 3.870 5.805 ;
        LAYER metal2 ;
        RECT  1.980 5.490 3.960 5.850 ;
        RECT  1.980 5.445 2.430 5.895 ;
        RECT  3.510 5.445 3.960 5.895 ;
    END
END or3_2

MACRO or3_1
    CLASS CORE ;
    FOREIGN or3_1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 5.490 1.800 5.850 ;
        END
    END ip2
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.005 2.160 4.365 3.420 ;
        RECT  2.835 5.490 4.230 5.850 ;
        RECT  3.870 3.060 4.230 5.850 ;
        RECT  3.465 7.110 3.825 9.270 ;
        RECT  2.835 7.110 3.825 7.470 ;
        RECT  2.835 5.490 3.195 7.470 ;
        END
    END op
    PIN ip3
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  3.060 4.680 3.420 5.040 ;
        END
    END ip3
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 4.680 0.990 5.040 ;
        END
    END ip1
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 5.670 0.990 ;
        RECT  3.195 0.000 3.555 2.790 ;
        RECT  1.575 0.000 1.935 2.790 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 5.670 11.340 ;
        RECT  2.610 8.010 2.970 11.340 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  0.765 2.160 1.125 3.780 ;
        RECT  2.385 2.160 2.745 3.780 ;
        RECT  0.765 3.420 2.745 3.780 ;
        RECT  2.025 6.255 2.475 6.705 ;
        RECT  2.070 3.420 2.430 7.470 ;
        RECT  0.765 7.110 2.430 7.470 ;
        RECT  0.765 7.110 1.125 9.270 ;
        RECT  3.510 6.255 3.960 6.705 ;
        LAYER via ;
        RECT  2.115 6.345 2.385 6.615 ;
        RECT  3.600 6.345 3.870 6.615 ;
        LAYER metal2 ;
        RECT  2.025 6.300 3.960 6.660 ;
        RECT  2.025 6.255 2.475 6.705 ;
        RECT  3.510 6.255 3.960 6.705 ;
    END
END or3_1

MACRO or2_4
    CLASS CORE ;
    FOREIGN or2_4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.860 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.060 2.160 3.420 9.270 ;
        END
    END op
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 4.680 1.800 5.040 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 3.870 0.990 4.230 ;
        END
    END ip1
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 4.860 11.340 ;
        RECT  3.825 6.750 4.185 11.340 ;
        RECT  2.250 6.750 2.610 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 4.860 0.990 ;
        RECT  3.870 0.000 4.230 3.420 ;
        RECT  2.250 0.000 2.610 3.420 ;
        RECT  0.630 0.000 0.990 3.420 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  1.440 2.160 1.800 4.230 ;
        RECT  1.440 3.870 2.610 4.230 ;
        RECT  2.250 3.870 2.610 5.670 ;
        RECT  0.855 5.310 2.745 5.670 ;
        RECT  0.855 5.310 1.215 9.270 ;
    END
END or2_4

MACRO or2_2
    CLASS CORE ;
    FOREIGN or2_2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.050 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 3.870 0.990 4.230 ;
        END
    END ip1
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 4.680 1.800 5.040 ;
        END
    END ip2
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.060 2.160 3.420 9.270 ;
        END
    END op
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 4.050 0.990 ;
        RECT  2.250 0.000 2.610 3.420 ;
        RECT  0.630 0.000 0.990 3.420 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 4.050 11.340 ;
        RECT  2.250 6.750 2.610 11.340 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  1.440 2.160 1.800 4.230 ;
        RECT  1.440 3.870 2.610 4.230 ;
        RECT  2.250 3.870 2.610 5.670 ;
        RECT  0.855 5.310 2.745 5.670 ;
        RECT  0.855 5.310 1.215 9.270 ;
    END
END or2_2

MACRO or2_1
    CLASS CORE ;
    FOREIGN or2_1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.050 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 3.870 0.990 4.230 ;
        END
    END ip1
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 4.680 1.800 5.040 ;
        END
    END ip2
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.060 2.160 3.420 9.270 ;
        END
    END op
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 4.050 0.990 ;
        RECT  2.250 0.000 2.610 2.790 ;
        RECT  0.630 0.000 0.990 2.790 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 4.050 11.340 ;
        RECT  2.250 8.010 2.610 11.340 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  1.440 2.160 1.800 4.230 ;
        RECT  1.440 3.870 2.610 4.230 ;
        RECT  2.250 3.870 2.610 5.670 ;
        RECT  0.855 5.310 2.745 5.670 ;
        RECT  0.855 5.310 1.215 9.270 ;
    END
END or2_1

MACRO not_ab_or_c_or_d
    CLASS CORE ;
    FOREIGN not_ab_or_c_or_d 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 3.870 0.990 4.230 ;
        END
    END ip1
    PIN ip3
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  3.060 5.490 3.420 5.850 ;
        END
    END ip3
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.680 5.490 5.040 9.270 ;
        RECT  3.870 5.490 5.040 5.850 ;
        RECT  3.870 2.160 4.230 5.850 ;
        RECT  2.250 3.060 4.230 3.420 ;
        RECT  2.250 2.160 2.610 3.420 ;
        END
    END op
    PIN ip4
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  4.680 3.870 5.040 4.230 ;
        END
    END ip4
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 4.680 2.610 5.040 ;
        END
    END ip2
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 5.670 11.340 ;
        RECT  2.250 8.010 2.610 11.340 ;
        RECT  0.630 8.010 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 5.670 0.990 ;
        RECT  4.680 0.000 5.040 2.790 ;
        RECT  3.060 0.000 3.420 2.790 ;
        RECT  0.630 0.000 0.990 2.790 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  1.440 7.110 3.420 7.470 ;
        RECT  1.440 7.110 1.800 9.270 ;
        RECT  3.060 7.110 3.420 9.270 ;
    END
END not_ab_or_c_or_d

MACRO nor4_4
    CLASS CORE ;
    FOREIGN nor4_4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.910 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 4.680 0.990 5.040 ;
        END
    END ip1
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.065 5.490 8.280 5.850 ;
        RECT  7.920 3.870 8.280 5.850 ;
        RECT  7.065 3.870 8.280 4.230 ;
        RECT  7.065 5.490 7.425 9.270 ;
        RECT  7.065 2.160 7.425 4.230 ;
        END
    END op
    PIN ip4
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  3.870 3.870 4.230 4.230 ;
        END
    END ip4
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 5.490 1.800 5.850 ;
        END
    END ip2
    PIN ip3
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 4.680 2.610 5.040 ;
        END
    END ip3
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 8.910 11.340 ;
        RECT  7.830 6.750 8.190 11.340 ;
        RECT  6.255 6.750 6.615 11.340 ;
        RECT  4.680 6.750 5.040 11.340 ;
        RECT  0.900 6.750 1.260 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 8.910 0.990 ;
        RECT  7.875 0.000 8.235 3.420 ;
        RECT  6.255 0.000 6.615 3.420 ;
        RECT  4.680 0.000 5.040 3.420 ;
        RECT  3.870 0.000 4.230 3.420 ;
        RECT  2.250 0.000 2.610 3.420 ;
        RECT  0.630 0.000 0.990 3.420 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  1.440 2.160 1.800 4.230 ;
        RECT  1.440 3.870 3.420 4.230 ;
        RECT  3.060 2.160 3.420 5.040 ;
        RECT  3.060 4.680 5.445 5.040 ;
        RECT  3.285 4.680 3.645 9.270 ;
        RECT  5.445 2.160 5.805 4.230 ;
        RECT  5.445 3.870 6.255 4.230 ;
        RECT  5.895 4.680 7.020 5.040 ;
        RECT  5.895 3.870 6.255 6.480 ;
        RECT  5.445 6.120 6.255 6.480 ;
        RECT  5.445 6.120 5.805 9.270 ;
    END
END nor4_4

MACRO nor4_2
    CLASS CORE ;
    FOREIGN nor4_2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.860 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip3
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 4.680 2.610 5.040 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 5.490 1.800 5.850 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 4.680 0.990 5.040 ;
        END
    END ip1
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.285 5.490 3.645 9.270 ;
        RECT  3.060 2.160 3.420 5.850 ;
        RECT  1.440 3.870 3.420 4.230 ;
        RECT  1.440 2.160 1.800 4.230 ;
        END
    END op
    PIN ip4
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  3.870 3.870 4.230 4.230 ;
        END
    END ip4
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 4.860 0.990 ;
        RECT  3.870 0.000 4.230 3.420 ;
        RECT  2.250 0.000 2.610 3.420 ;
        RECT  0.630 0.000 0.990 3.420 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 4.860 11.340 ;
        RECT  0.900 6.750 1.260 11.340 ;
        END
    END vdd!
END nor4_2

MACRO nor4_1
    CLASS CORE ;
    FOREIGN nor4_1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.860 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.285 5.490 3.645 9.270 ;
        RECT  3.060 2.160 3.420 5.850 ;
        RECT  1.440 3.060 3.420 3.420 ;
        RECT  1.440 2.160 1.800 3.420 ;
        END
    END op
    PIN ip4
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  3.870 3.870 4.230 4.230 ;
        END
    END ip4
    PIN ip3
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 4.680 2.610 5.040 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 5.490 1.800 5.850 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 6.300 0.990 6.660 ;
        END
    END ip1
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 4.860 0.990 ;
        RECT  3.870 0.000 4.230 2.790 ;
        RECT  2.250 0.000 2.610 2.790 ;
        RECT  0.630 0.000 0.990 2.790 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 4.860 11.340 ;
        RECT  0.900 8.010 1.260 11.340 ;
        END
    END vdd!
END nor4_1

MACRO nor3_4
    CLASS CORE ;
    FOREIGN nor3_4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.480 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.440 3.870 4.995 4.230 ;
        RECT  4.635 2.160 4.995 4.230 ;
        RECT  3.060 2.160 3.420 5.850 ;
        RECT  2.970 5.490 3.330 9.270 ;
        RECT  1.440 2.160 1.800 4.230 ;
        END
    END op
    PIN ip3
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 4.680 2.610 5.040 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  4.140 5.535 4.410 5.805 ;
        RECT  1.485 5.535 1.755 5.805 ;
        LAYER metal2 ;
        RECT  4.050 5.445 4.500 5.895 ;
        RECT  1.395 5.490 4.500 5.850 ;
        RECT  1.395 5.445 1.845 5.895 ;
        LAYER metal1 ;
        RECT  4.050 5.445 4.500 5.895 ;
        RECT  1.395 5.445 1.845 5.895 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  5.085 6.345 5.355 6.615 ;
        RECT  0.720 6.345 0.990 6.615 ;
        LAYER metal2 ;
        RECT  4.995 6.255 5.445 6.705 ;
        RECT  0.630 6.300 5.445 6.660 ;
        RECT  0.630 6.255 1.080 6.705 ;
        LAYER metal1 ;
        RECT  4.995 6.255 5.445 6.705 ;
        RECT  0.630 6.255 1.080 6.705 ;
        END
    END ip1
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 6.480 11.340 ;
        RECT  4.860 6.975 5.220 11.340 ;
        RECT  1.125 6.975 1.485 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 6.480 0.990 ;
        RECT  5.445 0.000 5.805 3.420 ;
        RECT  3.825 0.000 4.185 3.420 ;
        RECT  2.295 0.000 2.655 3.420 ;
        RECT  0.630 0.000 0.990 3.420 ;
        END
    END gnd!
END nor3_4

MACRO nor3_2
    CLASS CORE ;
    FOREIGN nor3_2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.050 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.060 3.870 3.420 5.850 ;
        RECT  2.790 5.490 3.150 9.270 ;
        RECT  1.350 3.870 3.420 4.230 ;
        RECT  2.790 2.160 3.150 4.230 ;
        RECT  1.350 2.160 1.710 4.230 ;
        END
    END op
    PIN ip3
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 4.680 2.610 5.040 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 5.490 1.800 5.850 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 3.870 0.990 4.230 ;
        END
    END ip1
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 4.050 0.990 ;
        RECT  2.070 0.000 2.430 3.420 ;
        RECT  0.630 0.000 0.990 3.420 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 4.050 11.340 ;
        RECT  0.900 6.750 1.260 11.340 ;
        END
    END vdd!
END nor3_2

MACRO nor3_1
    CLASS CORE ;
    FOREIGN nor3_1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.050 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.060 3.870 3.420 5.850 ;
        RECT  2.790 5.490 3.150 9.270 ;
        RECT  1.350 3.870 3.420 4.230 ;
        RECT  2.790 2.160 3.150 4.230 ;
        RECT  1.350 2.160 1.710 4.230 ;
        END
    END op
    PIN ip3
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 4.680 2.610 5.040 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 5.490 1.800 5.850 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 6.345 0.990 6.705 ;
        END
    END ip1
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 4.050 0.990 ;
        RECT  2.070 0.000 2.430 2.790 ;
        RECT  0.630 0.000 0.990 2.790 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 4.050 11.340 ;
        RECT  0.900 8.010 1.260 11.340 ;
        END
    END vdd!
END nor3_1

MACRO nor2_4
    CLASS CORE ;
    FOREIGN nor2_4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  3.105 5.535 3.375 5.805 ;
        RECT  0.720 5.535 0.990 5.805 ;
        LAYER metal2 ;
        RECT  3.015 5.445 3.465 5.895 ;
        RECT  0.630 5.490 3.465 5.850 ;
        RECT  0.630 5.445 1.080 5.895 ;
        LAYER metal1 ;
        RECT  3.015 5.445 3.465 5.895 ;
        RECT  0.630 5.445 1.080 5.895 ;
        END
    END ip1
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  3.915 4.725 4.185 4.995 ;
        RECT  1.485 4.725 1.755 4.995 ;
        LAYER metal2 ;
        RECT  3.825 4.635 4.275 5.085 ;
        RECT  1.395 4.680 4.275 5.040 ;
        RECT  1.395 4.635 1.845 5.085 ;
        LAYER metal1 ;
        RECT  3.825 4.635 4.275 5.085 ;
        RECT  1.395 4.635 1.845 5.085 ;
        END
    END ip2
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.680 3.870 5.040 9.270 ;
        RECT  1.440 3.870 5.040 4.230 ;
        RECT  3.870 2.160 4.230 4.230 ;
        RECT  2.250 3.870 2.610 9.270 ;
        RECT  1.440 2.160 1.800 4.230 ;
        END
    END op
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 5.670 11.340 ;
        RECT  3.330 6.750 3.690 11.340 ;
        RECT  0.900 6.750 1.260 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 5.670 0.990 ;
        RECT  4.680 0.000 5.040 3.420 ;
        RECT  3.060 0.000 3.420 3.420 ;
        RECT  2.250 0.000 2.610 3.420 ;
        RECT  0.630 0.000 0.990 3.420 ;
        END
    END gnd!
END nor2_4

MACRO nor2_2
    CLASS CORE ;
    FOREIGN nor2_2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.240 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.250 3.870 2.610 9.270 ;
        RECT  1.440 3.870 2.610 4.230 ;
        RECT  1.440 2.160 1.800 4.230 ;
        END
    END op
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 4.680 1.800 5.040 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip1
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 3.240 0.990 ;
        RECT  2.250 0.000 2.610 3.420 ;
        RECT  0.630 0.000 0.990 3.420 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 3.240 11.340 ;
        RECT  0.900 6.750 1.260 11.340 ;
        END
    END vdd!
END nor2_2

MACRO nor2_1
    CLASS CORE ;
    FOREIGN nor2_1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.240 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.250 3.870 2.610 9.270 ;
        RECT  1.440 3.870 2.610 4.230 ;
        RECT  1.440 2.160 1.800 4.230 ;
        END
    END op
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 4.680 1.800 5.040 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip1
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 3.240 0.990 ;
        RECT  2.250 0.000 2.610 2.790 ;
        RECT  0.630 0.000 0.990 2.790 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 3.240 11.340 ;
        RECT  0.900 8.010 1.260 11.340 ;
        END
    END vdd!
END nor2_1

MACRO nand4_4
    CLASS CORE ;
    FOREIGN nand4_4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.100 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 3.870 2.610 4.230 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip1
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.300 5.490 7.470 5.850 ;
        RECT  7.110 3.870 7.470 5.850 ;
        RECT  6.300 3.870 7.470 4.230 ;
        RECT  6.300 5.490 6.660 9.270 ;
        RECT  6.300 2.160 6.660 4.230 ;
        END
    END op
    PIN ip3
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 4.680 2.610 5.040 ;
        END
    END ip3
    PIN ip4
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  3.870 4.680 4.230 5.040 ;
        END
    END ip4
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 8.100 11.340 ;
        RECT  7.110 6.750 7.470 11.340 ;
        RECT  5.490 7.290 5.850 11.340 ;
        RECT  3.870 6.750 4.230 11.340 ;
        RECT  2.250 6.750 2.610 11.340 ;
        RECT  0.630 6.750 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 8.100 0.990 ;
        RECT  7.110 0.000 7.470 3.420 ;
        RECT  5.490 0.000 5.850 3.420 ;
        RECT  3.870 0.000 4.230 3.420 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  0.630 2.160 0.990 5.040 ;
        RECT  0.630 4.680 1.800 5.040 ;
        RECT  1.440 5.490 4.635 5.850 ;
        RECT  1.440 4.680 1.800 9.270 ;
        RECT  3.060 5.490 3.420 9.270 ;
        RECT  4.680 2.160 5.040 4.230 ;
        RECT  4.680 3.870 5.490 4.230 ;
        RECT  5.130 4.680 6.255 5.040 ;
        RECT  5.130 3.870 5.490 6.660 ;
        RECT  4.680 6.300 5.490 6.660 ;
        RECT  4.680 6.300 5.040 9.270 ;
    END
END nand4_4

MACRO nand4_2
    CLASS CORE ;
    FOREIGN nand4_2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.860 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.250 4.680 4.230 5.040 ;
        RECT  3.870 2.160 4.230 5.040 ;
        RECT  3.060 6.030 3.420 9.270 ;
        RECT  1.440 6.030 3.420 6.390 ;
        RECT  2.250 4.680 2.610 6.390 ;
        RECT  1.440 6.030 1.800 9.270 ;
        END
    END op
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip1
    PIN ip4
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  3.870 5.490 4.230 5.850 ;
        END
    END ip4
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 4.680 1.800 5.040 ;
        END
    END ip2
    PIN ip3
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 3.870 2.610 4.230 ;
        END
    END ip3
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 4.860 11.340 ;
        RECT  3.870 6.750 4.230 11.340 ;
        RECT  2.250 6.750 2.610 11.340 ;
        RECT  0.630 6.750 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 4.860 0.990 ;
        RECT  0.630 0.000 0.990 3.420 ;
        END
    END gnd!
END nand4_2

MACRO nand4_1
    CLASS CORE ;
    FOREIGN nand4_1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.860 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip4
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  3.870 6.300 4.230 6.660 ;
        END
    END ip4
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 4.680 1.800 5.040 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip1
    PIN ip3
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 3.060 2.610 3.420 ;
        END
    END ip3
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.250 5.490 4.230 5.850 ;
        RECT  3.870 2.160 4.230 5.850 ;
        RECT  3.060 7.110 3.420 9.270 ;
        RECT  1.440 7.110 3.420 7.470 ;
        RECT  2.250 5.490 2.610 7.470 ;
        RECT  1.440 7.110 1.800 9.270 ;
        END
    END op
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 4.860 11.340 ;
        RECT  3.870 8.010 4.230 11.340 ;
        RECT  2.250 8.010 2.610 11.340 ;
        RECT  0.630 8.010 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 4.860 0.990 ;
        RECT  0.630 0.000 0.990 2.790 ;
        END
    END gnd!
END nand4_1

MACRO nand3_4
    CLASS CORE ;
    FOREIGN nand3_4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.480 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  5.535 5.535 5.805 5.805 ;
        RECT  0.675 5.535 0.945 5.805 ;
        LAYER metal2 ;
        RECT  5.445 5.445 5.895 5.895 ;
        RECT  0.585 5.490 5.895 5.850 ;
        RECT  0.585 5.445 1.035 5.895 ;
        LAYER metal1 ;
        RECT  5.445 5.445 5.895 5.895 ;
        RECT  0.585 5.445 1.035 5.895 ;
        END
    END ip1
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  3.915 4.725 4.185 4.995 ;
        RECT  1.485 4.725 1.755 4.995 ;
        LAYER metal2 ;
        RECT  3.825 4.635 4.275 5.085 ;
        RECT  1.395 4.680 4.275 5.040 ;
        RECT  1.395 4.635 1.845 5.085 ;
        LAYER metal1 ;
        RECT  3.825 4.635 4.275 5.085 ;
        RECT  1.395 4.635 1.845 5.085 ;
        END
    END ip2
    PIN ip3
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  3.060 3.870 3.420 4.230 ;
        END
    END ip3
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.310 6.300 5.670 9.270 ;
        RECT  3.735 6.300 5.670 6.660 ;
        RECT  4.500 5.490 4.860 6.660 ;
        RECT  1.440 5.490 4.860 5.850 ;
        RECT  3.735 6.300 4.095 9.270 ;
        RECT  2.250 3.240 3.105 3.600 ;
        RECT  2.745 2.160 3.105 3.600 ;
        RECT  2.250 3.240 2.610 5.850 ;
        RECT  2.205 6.300 2.565 9.270 ;
        RECT  0.630 6.300 2.565 6.660 ;
        RECT  1.440 5.490 1.800 6.660 ;
        RECT  0.630 6.300 0.990 9.270 ;
        END
    END op
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 6.480 11.340 ;
        RECT  4.545 6.930 4.905 11.340 ;
        RECT  2.970 6.750 3.330 11.340 ;
        RECT  1.395 6.930 1.755 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 6.480 0.990 ;
        RECT  4.590 0.000 4.950 3.420 ;
        RECT  0.900 0.000 1.260 3.420 ;
        END
    END gnd!
END nand3_4

MACRO nand3_2
    CLASS CORE ;
    FOREIGN nand3_2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.050 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.250 3.240 3.105 3.600 ;
        RECT  2.745 2.160 3.105 3.600 ;
        RECT  1.440 5.490 2.610 5.850 ;
        RECT  2.250 3.240 2.610 5.850 ;
        RECT  2.205 6.300 2.565 9.270 ;
        RECT  0.630 6.300 2.565 6.660 ;
        RECT  1.440 5.490 1.800 6.660 ;
        RECT  0.630 6.300 0.990 9.270 ;
        END
    END op
    PIN ip3
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  3.060 3.870 3.420 4.230 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 4.680 1.800 5.040 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  0.675 5.535 0.945 5.805 ;
        LAYER metal2 ;
        RECT  0.585 5.445 1.035 5.895 ;
        LAYER metal1 ;
        RECT  0.585 5.445 1.035 5.895 ;
        END
    END ip1
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 4.050 0.990 ;
        RECT  0.900 0.000 1.260 3.420 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 4.050 11.340 ;
        RECT  2.970 6.750 3.330 11.340 ;
        RECT  1.395 6.930 1.755 11.340 ;
        END
    END vdd!
END nand3_2

MACRO nand3_1
    CLASS CORE ;
    FOREIGN nand3_1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.050 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip3
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  3.060 3.870 3.420 4.230 ;
        END
    END ip3
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.970 6.300 3.330 9.270 ;
        RECT  2.250 2.250 3.105 2.610 ;
        RECT  1.395 6.300 3.330 6.660 ;
        RECT  2.250 2.250 2.610 6.660 ;
        RECT  1.395 6.300 1.755 9.270 ;
        END
    END op
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 4.680 1.800 5.040 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  0.675 5.535 0.945 5.805 ;
        LAYER metal2 ;
        RECT  0.585 5.445 1.035 5.895 ;
        LAYER metal1 ;
        RECT  0.585 5.445 1.035 5.895 ;
        END
    END ip1
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 4.050 0.990 ;
        RECT  0.900 0.000 1.260 2.790 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 4.050 11.340 ;
        RECT  2.205 8.010 2.565 11.340 ;
        RECT  0.630 8.010 0.990 11.340 ;
        END
    END vdd!
END nand3_1

MACRO nand2_4
    CLASS CORE ;
    FOREIGN nand2_4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.860 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  3.870 5.535 4.140 5.805 ;
        RECT  0.720 5.535 0.990 5.805 ;
        LAYER metal2 ;
        RECT  3.780 5.445 4.230 5.895 ;
        RECT  0.630 5.490 4.230 5.850 ;
        RECT  0.630 5.445 1.080 5.895 ;
        LAYER metal1 ;
        RECT  3.780 5.445 4.230 5.895 ;
        RECT  0.630 5.445 1.080 5.895 ;
        END
    END ip1
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 4.680 1.800 5.040 ;
        END
    END ip2
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.970 6.300 3.330 9.270 ;
        RECT  1.440 6.300 3.330 6.660 ;
        RECT  2.250 2.160 2.610 6.660 ;
        RECT  1.440 6.300 1.800 9.270 ;
        END
    END op
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 4.860 0.990 ;
        RECT  3.690 0.000 4.050 3.420 ;
        RECT  0.945 0.000 1.305 3.420 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 4.860 11.340 ;
        RECT  3.780 7.065 4.140 11.340 ;
        RECT  2.205 7.065 2.565 11.340 ;
        RECT  0.630 7.065 0.990 11.340 ;
        END
    END vdd!
END nand2_4

MACRO nand2_2
    CLASS CORE ;
    FOREIGN nand2_2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.240 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip1
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 4.680 1.800 5.040 ;
        END
    END ip2
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.440 6.300 2.610 6.660 ;
        RECT  2.250 2.160 2.610 6.660 ;
        RECT  1.440 6.300 1.800 9.270 ;
        END
    END op
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 3.240 0.990 ;
        RECT  0.945 0.000 1.305 3.420 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 3.240 11.340 ;
        RECT  2.205 7.065 2.565 11.340 ;
        RECT  0.630 6.750 0.990 11.340 ;
        END
    END vdd!
END nand2_2

MACRO nand2_1
    CLASS CORE ;
    FOREIGN nand2_1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.240 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip1
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 4.680 1.800 5.040 ;
        END
    END ip2
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.440 7.245 2.610 7.605 ;
        RECT  2.250 2.160 2.610 7.605 ;
        RECT  1.440 7.245 1.800 9.270 ;
        END
    END op
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 3.240 0.990 ;
        RECT  0.945 0.000 1.305 2.655 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 3.240 11.340 ;
        RECT  2.205 8.055 2.565 11.340 ;
        RECT  0.630 8.055 0.990 11.340 ;
        END
    END vdd!
END nand2_1

MACRO mux4_2
    CLASS CORE ;
    FOREIGN mux4_2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.250 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN s1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  10.710 4.725 10.980 4.995 ;
        RECT  7.965 4.725 8.235 4.995 ;
        LAYER metal2 ;
        RECT  10.620 4.635 11.070 5.085 ;
        RECT  7.875 4.680 11.070 5.040 ;
        RECT  7.875 4.635 8.325 5.085 ;
        LAYER metal1 ;
        RECT  10.620 4.635 11.070 5.085 ;
        RECT  7.875 4.635 8.325 5.085 ;
        END
    END s1
    PIN s0
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  15.660 5.535 15.930 5.805 ;
        RECT  14.040 5.535 14.310 5.805 ;
        RECT  4.995 5.535 5.265 5.805 ;
        RECT  1.485 5.535 1.755 5.805 ;
        LAYER metal2 ;
        RECT  15.570 5.445 16.020 5.895 ;
        RECT  1.395 5.490 16.020 5.850 ;
        RECT  13.950 5.445 14.400 5.895 ;
        RECT  4.905 5.445 5.355 5.895 ;
        RECT  1.395 5.445 1.845 5.895 ;
        LAYER metal1 ;
        RECT  15.570 5.445 16.020 5.895 ;
        RECT  13.950 5.445 14.400 5.895 ;
        RECT  4.905 5.445 5.355 5.895 ;
        RECT  1.395 5.445 1.845 5.895 ;
        END
    END s0
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  6.300 4.680 6.660 5.040 ;
        END
    END ip2
    PIN ip3
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  11.970 4.680 12.330 5.040 ;
        END
    END ip3
    PIN ip4
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  16.830 3.870 17.190 4.230 ;
        END
    END ip4
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  18.045 6.300 18.810 6.660 ;
        RECT  18.450 3.870 18.810 6.660 ;
        RECT  18.045 3.870 18.810 4.230 ;
        RECT  18.045 6.300 18.405 9.270 ;
        RECT  18.045 2.160 18.405 4.230 ;
        END
    END op
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 4.680 0.990 5.040 ;
        END
    END ip1
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 20.250 0.990 ;
        RECT  17.235 0.000 17.595 3.420 ;
        RECT  11.970 0.000 12.330 3.420 ;
        RECT  7.110 0.000 7.470 3.420 ;
        RECT  1.440 0.000 1.800 3.420 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 20.250 11.340 ;
        RECT  17.235 6.750 17.595 11.340 ;
        RECT  11.970 6.750 12.330 11.340 ;
        RECT  7.110 6.750 7.470 11.340 ;
        RECT  1.395 6.750 1.755 11.340 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  0.630 8.685 1.080 9.135 ;
        RECT  0.630 6.750 0.990 9.270 ;
        RECT  0.630 2.205 1.080 2.655 ;
        RECT  0.630 2.160 0.990 3.420 ;
        RECT  2.250 3.825 2.880 4.275 ;
        RECT  2.250 2.160 2.610 9.270 ;
        RECT  3.330 2.205 3.780 2.655 ;
        RECT  3.375 8.685 3.825 9.135 ;
        RECT  3.375 2.160 3.735 9.270 ;
        RECT  4.140 6.255 4.590 6.705 ;
        RECT  4.185 2.160 4.545 9.270 ;
        RECT  4.995 2.160 5.355 4.230 ;
        RECT  6.300 2.160 6.660 4.230 ;
        RECT  4.995 3.870 6.660 4.230 ;
        RECT  5.670 3.870 6.030 8.370 ;
        RECT  4.995 8.010 6.660 8.370 ;
        RECT  4.995 8.010 5.355 9.270 ;
        RECT  6.300 6.750 6.660 9.270 ;
        RECT  7.920 2.160 8.280 4.230 ;
        RECT  7.110 3.870 8.640 4.230 ;
        RECT  7.110 3.870 7.470 6.300 ;
        RECT  7.110 5.940 8.280 6.300 ;
        RECT  7.920 5.940 8.280 9.270 ;
        RECT  9.090 6.255 9.540 6.705 ;
        RECT  9.135 2.160 9.495 9.270 ;
        RECT  9.900 7.065 10.350 7.515 ;
        RECT  9.945 2.160 10.305 9.270 ;
        RECT  10.755 2.160 11.115 4.275 ;
        RECT  10.755 3.915 11.700 4.275 ;
        RECT  11.340 3.915 11.700 5.805 ;
        RECT  10.755 5.445 11.700 5.805 ;
        RECT  10.710 6.255 11.160 6.705 ;
        RECT  10.755 5.445 11.115 9.270 ;
        RECT  12.780 2.250 14.355 2.610 ;
        RECT  13.995 2.160 14.355 2.790 ;
        RECT  12.780 2.160 13.140 9.270 ;
        RECT  13.590 8.010 13.950 9.270 ;
        RECT  12.780 8.910 13.950 9.270 ;
        RECT  13.950 3.825 14.400 4.275 ;
        RECT  14.715 6.255 15.165 6.705 ;
        RECT  14.760 2.160 15.120 6.795 ;
        RECT  14.400 6.435 14.760 9.270 ;
        RECT  15.615 2.250 16.785 2.610 ;
        RECT  16.425 2.160 16.785 3.420 ;
        RECT  15.615 2.160 15.975 5.085 ;
        RECT  15.615 4.725 16.785 5.085 ;
        RECT  15.210 8.010 15.570 9.270 ;
        RECT  16.425 4.725 16.785 9.270 ;
        RECT  15.210 8.910 16.785 9.270 ;
        RECT  17.595 5.445 18.045 5.895 ;
        LAYER via ;
        RECT  0.720 8.775 0.990 9.045 ;
        RECT  0.720 2.295 0.990 2.565 ;
        RECT  2.520 3.915 2.790 4.185 ;
        RECT  3.420 2.295 3.690 2.565 ;
        RECT  3.465 8.775 3.735 9.045 ;
        RECT  4.230 6.345 4.500 6.615 ;
        RECT  9.180 6.345 9.450 6.615 ;
        RECT  9.990 7.155 10.260 7.425 ;
        RECT  10.800 6.345 11.070 6.615 ;
        RECT  14.040 3.915 14.310 4.185 ;
        RECT  14.805 6.345 15.075 6.615 ;
        RECT  17.685 5.535 17.955 5.805 ;
        LAYER metal2 ;
        RECT  0.630 2.250 3.780 2.610 ;
        RECT  0.630 2.205 1.080 2.655 ;
        RECT  3.330 2.205 3.780 2.655 ;
        RECT  0.630 8.730 3.825 9.090 ;
        RECT  0.630 8.685 1.080 9.135 ;
        RECT  3.375 8.685 3.825 9.135 ;
        RECT  4.140 6.300 9.540 6.660 ;
        RECT  4.140 6.255 4.590 6.705 ;
        RECT  9.090 6.255 9.540 6.705 ;
        RECT  2.430 3.870 14.400 4.230 ;
        RECT  2.430 3.825 2.880 4.275 ;
        RECT  13.950 3.825 14.400 4.275 ;
        RECT  10.710 6.300 15.165 6.660 ;
        RECT  10.710 6.255 11.160 6.705 ;
        RECT  14.715 6.255 15.165 6.705 ;
        RECT  17.595 5.445 18.045 5.895 ;
        RECT  17.640 5.445 18.000 7.470 ;
        RECT  9.900 7.110 18.000 7.470 ;
        RECT  9.900 7.065 10.350 7.515 ;
    END
END mux4_2

MACRO mux3_2
    CLASS CORE ;
    FOREIGN mux3_2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.390 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 4.680 0.990 5.040 ;
        END
    END ip1
    PIN s0
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  4.995 5.535 5.265 5.805 ;
        RECT  1.485 5.535 1.755 5.805 ;
        LAYER metal2 ;
        RECT  4.905 5.445 5.355 5.895 ;
        RECT  1.395 5.490 5.355 5.850 ;
        RECT  1.395 5.445 1.845 5.895 ;
        LAYER metal1 ;
        RECT  4.905 5.445 5.355 5.895 ;
        RECT  1.395 5.445 1.845 5.895 ;
        END
    END s0
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  6.300 5.490 6.660 5.850 ;
        END
    END ip2
    PIN s1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  10.845 4.725 11.115 4.995 ;
        RECT  7.965 4.725 8.235 4.995 ;
        LAYER metal2 ;
        RECT  10.755 4.635 11.205 5.085 ;
        RECT  7.875 4.680 11.205 5.040 ;
        RECT  7.875 4.635 8.325 5.085 ;
        LAYER metal1 ;
        RECT  10.755 4.635 11.205 5.085 ;
        RECT  7.875 4.635 8.325 5.085 ;
        END
    END s1
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.770 6.300 14.760 6.660 ;
        RECT  14.400 3.870 14.760 6.660 ;
        RECT  13.770 3.870 14.760 4.230 ;
        RECT  13.770 6.300 14.130 9.270 ;
        RECT  13.770 2.160 14.130 4.230 ;
        END
    END op
    PIN ip3
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  12.780 4.680 13.140 5.040 ;
        END
    END ip3
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 15.390 11.340 ;
        RECT  12.960 6.750 13.320 11.340 ;
        RECT  7.110 6.750 7.470 11.340 ;
        RECT  1.440 6.750 1.800 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 15.390 0.990 ;
        RECT  12.960 0.000 13.320 3.420 ;
        RECT  7.110 0.000 7.470 3.420 ;
        RECT  1.440 0.000 1.800 3.420 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  0.630 8.685 1.080 9.135 ;
        RECT  0.630 6.750 0.990 9.270 ;
        RECT  0.630 2.205 1.080 2.655 ;
        RECT  0.630 2.160 0.990 3.420 ;
        RECT  2.250 3.870 2.880 4.230 ;
        RECT  2.250 2.160 2.610 9.270 ;
        RECT  3.330 2.205 3.780 2.655 ;
        RECT  3.330 8.685 3.780 9.135 ;
        RECT  3.375 2.160 3.735 9.270 ;
        RECT  4.140 6.255 4.590 6.705 ;
        RECT  4.185 2.160 4.545 9.270 ;
        RECT  4.995 2.160 5.355 4.230 ;
        RECT  6.300 2.160 6.660 4.230 ;
        RECT  4.995 3.870 6.660 4.230 ;
        RECT  5.670 3.870 6.030 6.660 ;
        RECT  4.995 6.300 6.660 6.660 ;
        RECT  4.995 6.300 5.355 9.270 ;
        RECT  6.300 6.300 6.660 9.270 ;
        RECT  7.920 2.160 8.280 4.230 ;
        RECT  7.920 3.870 8.955 4.230 ;
        RECT  8.595 3.870 8.955 5.850 ;
        RECT  7.920 5.490 8.955 5.850 ;
        RECT  7.920 5.490 8.280 9.270 ;
        RECT  9.180 6.255 9.630 6.705 ;
        RECT  9.225 2.160 9.585 9.270 ;
        RECT  9.990 5.445 10.440 5.895 ;
        RECT  10.035 2.160 10.395 9.270 ;
        RECT  10.845 2.250 12.510 2.610 ;
        RECT  12.150 2.160 12.510 3.420 ;
        RECT  10.845 2.160 11.205 4.230 ;
        RECT  10.845 3.870 11.880 4.230 ;
        RECT  11.520 3.870 11.880 6.660 ;
        RECT  10.845 6.300 11.880 6.660 ;
        RECT  10.845 6.300 11.205 9.270 ;
        RECT  12.150 6.750 12.510 9.270 ;
        RECT  10.845 8.910 12.510 9.270 ;
        RECT  13.320 5.445 13.770 5.895 ;
        LAYER via ;
        RECT  0.720 8.775 0.990 9.045 ;
        RECT  0.720 2.295 0.990 2.565 ;
        RECT  3.420 8.775 3.690 9.045 ;
        RECT  3.420 2.295 3.690 2.565 ;
        RECT  4.230 6.345 4.500 6.615 ;
        RECT  9.270 6.345 9.540 6.615 ;
        RECT  10.080 5.535 10.350 5.805 ;
        RECT  13.410 5.535 13.680 5.805 ;
        LAYER metal2 ;
        RECT  0.630 8.730 3.780 9.090 ;
        RECT  0.630 8.685 1.080 9.135 ;
        RECT  3.330 8.685 3.780 9.135 ;
        RECT  0.630 2.250 3.780 2.610 ;
        RECT  0.630 2.205 1.080 2.655 ;
        RECT  3.330 2.205 3.780 2.655 ;
        RECT  4.140 6.300 9.630 6.660 ;
        RECT  4.140 6.255 4.590 6.705 ;
        RECT  9.180 6.255 9.630 6.705 ;
        RECT  9.990 5.490 13.770 5.850 ;
        RECT  9.990 5.445 10.440 5.895 ;
        RECT  13.320 5.445 13.770 5.895 ;
    END
END mux3_2

MACRO mux2_4
    CLASS CORE ;
    FOREIGN mux2_4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.290 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.490 2.160 5.850 9.270 ;
        END
    END op
    PIN s
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  3.915 6.345 4.185 6.615 ;
        RECT  1.485 6.345 1.755 6.615 ;
        LAYER metal2 ;
        RECT  3.825 6.255 4.275 6.705 ;
        RECT  1.395 6.300 4.275 6.660 ;
        RECT  1.395 6.255 1.845 6.705 ;
        LAYER metal1 ;
        RECT  3.825 6.255 4.275 6.705 ;
        RECT  1.395 6.255 1.845 6.705 ;
        END
    END s
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  3.870 5.490 4.230 5.850 ;
        END
    END ip1
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 4.680 2.610 5.040 ;
        END
    END ip2
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 7.290 11.340 ;
        RECT  6.210 6.750 6.570 11.340 ;
        RECT  4.770 6.750 5.130 11.340 ;
        RECT  3.915 8.010 4.275 11.340 ;
        RECT  1.350 8.010 1.710 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 7.290 0.990 ;
        RECT  6.210 0.000 6.570 3.420 ;
        RECT  4.770 0.000 5.130 3.420 ;
        RECT  3.915 0.000 4.275 2.790 ;
        RECT  1.350 0.000 1.710 2.790 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  0.630 3.870 1.845 4.230 ;
        RECT  1.395 3.825 1.845 4.275 ;
        RECT  0.630 2.160 0.990 9.270 ;
        RECT  3.825 3.825 4.275 4.275 ;
        RECT  2.655 2.160 3.015 3.420 ;
        RECT  2.655 3.060 3.420 3.420 ;
        RECT  3.060 4.680 5.040 5.040 ;
        RECT  3.060 3.060 3.420 5.850 ;
        RECT  2.655 5.490 3.420 5.850 ;
        RECT  2.655 5.490 3.015 9.270 ;
        LAYER via ;
        RECT  1.485 3.915 1.755 4.185 ;
        RECT  3.915 3.915 4.185 4.185 ;
        LAYER metal2 ;
        RECT  1.395 3.870 4.275 4.230 ;
        RECT  1.395 3.825 1.845 4.275 ;
        RECT  3.825 3.825 4.275 4.275 ;
    END
END mux2_4

MACRO mux2_2
    CLASS CORE ;
    FOREIGN mux2_2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.480 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 4.680 2.610 5.040 ;
        END
    END ip2
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.490 2.160 5.850 9.270 ;
        END
    END op
    PIN s
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  3.915 6.345 4.185 6.615 ;
        RECT  1.485 6.345 1.755 6.615 ;
        LAYER metal2 ;
        RECT  3.825 6.255 4.275 6.705 ;
        RECT  1.395 6.300 4.275 6.660 ;
        RECT  1.395 6.255 1.845 6.705 ;
        LAYER metal1 ;
        RECT  3.825 6.255 4.275 6.705 ;
        RECT  1.395 6.255 1.845 6.705 ;
        END
    END s
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  3.825 5.580 4.230 5.850 ;
        RECT  3.870 5.490 4.230 5.850 ;
        END
    END ip1
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 6.480 11.340 ;
        RECT  4.770 6.750 5.130 11.340 ;
        RECT  3.915 8.010 4.275 11.340 ;
        RECT  1.350 8.010 1.710 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 6.480 0.990 ;
        RECT  4.770 0.000 5.130 3.420 ;
        RECT  3.915 0.000 4.275 2.790 ;
        RECT  1.350 0.000 1.710 2.790 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  0.630 3.870 1.845 4.230 ;
        RECT  1.395 3.825 1.845 4.275 ;
        RECT  0.630 2.160 0.990 9.270 ;
        RECT  3.825 3.825 4.275 4.275 ;
        RECT  2.655 2.160 3.015 3.420 ;
        RECT  2.655 3.060 3.420 3.420 ;
        RECT  3.060 4.680 5.040 5.040 ;
        RECT  3.060 3.060 3.420 5.850 ;
        RECT  2.655 5.490 3.420 5.850 ;
        RECT  2.655 5.490 3.015 9.270 ;
        LAYER via ;
        RECT  1.485 3.915 1.755 4.185 ;
        RECT  3.915 3.915 4.185 4.185 ;
        LAYER metal2 ;
        RECT  1.395 3.870 4.275 4.230 ;
        RECT  1.395 3.825 1.845 4.275 ;
        RECT  3.825 3.825 4.275 4.275 ;
    END
END mux2_2

MACRO mux2_1
    CLASS CORE ;
    FOREIGN mux2_1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.480 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.490 2.160 5.850 9.270 ;
        END
    END op
    PIN s
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  3.915 6.345 4.185 6.615 ;
        RECT  1.485 6.345 1.755 6.615 ;
        LAYER metal2 ;
        RECT  3.825 6.255 4.275 6.705 ;
        RECT  1.395 6.300 4.275 6.660 ;
        RECT  1.395 6.255 1.845 6.705 ;
        LAYER metal1 ;
        RECT  3.825 6.255 4.275 6.705 ;
        RECT  1.395 6.255 1.845 6.705 ;
        END
    END s
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  3.870 5.490 4.230 5.850 ;
        END
    END ip1
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 4.680 2.610 5.040 ;
        END
    END ip2
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 6.480 11.340 ;
        RECT  4.770 8.010 5.130 11.340 ;
        RECT  3.915 8.010 4.275 11.340 ;
        RECT  1.350 8.010 1.710 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 6.480 0.990 ;
        RECT  4.770 0.000 5.130 2.790 ;
        RECT  3.915 0.000 4.275 2.790 ;
        RECT  1.350 0.000 1.710 2.790 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  0.630 3.870 1.845 4.230 ;
        RECT  1.395 3.825 1.845 4.275 ;
        RECT  0.630 2.160 0.990 9.270 ;
        RECT  3.825 3.825 4.275 4.275 ;
        RECT  2.655 2.160 3.015 3.420 ;
        RECT  2.655 3.060 3.420 3.420 ;
        RECT  3.060 4.680 5.040 5.040 ;
        RECT  3.060 3.060 3.420 5.850 ;
        RECT  2.655 5.490 3.420 5.850 ;
        RECT  2.655 5.490 3.015 9.270 ;
        LAYER via ;
        RECT  1.485 3.915 1.755 4.185 ;
        RECT  3.915 3.915 4.185 4.185 ;
        LAYER metal2 ;
        RECT  1.395 3.870 4.275 4.230 ;
        RECT  1.395 3.825 1.845 4.275 ;
        RECT  3.825 3.825 4.275 4.275 ;
    END
END mux2_1

MACRO lrsp_4
    CLASS CORE ;
    FOREIGN lrsp_4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.770 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN s
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  7.155 3.915 7.425 4.185 ;
        RECT  1.485 3.915 1.755 4.185 ;
        LAYER metal2 ;
        RECT  7.065 3.825 7.515 4.275 ;
        RECT  1.395 3.870 7.515 4.230 ;
        RECT  1.395 3.825 1.845 4.275 ;
        LAYER metal1 ;
        RECT  7.065 3.825 7.515 4.275 ;
        RECT  1.395 3.825 1.845 4.275 ;
        END
    END s
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.610 5.490 11.970 9.270 ;
        RECT  11.160 3.870 11.970 4.230 ;
        RECT  11.610 2.160 11.970 4.230 ;
        RECT  11.160 5.490 11.970 5.850 ;
        RECT  11.160 3.870 11.520 5.850 ;
        RECT  7.920 4.680 11.520 5.040 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  8.775 6.345 9.045 6.615 ;
        RECT  2.295 6.345 2.565 6.615 ;
        LAYER metal2 ;
        RECT  8.685 6.255 9.135 6.705 ;
        RECT  2.205 6.300 9.135 6.660 ;
        RECT  2.205 6.255 2.655 6.705 ;
        LAYER metal1 ;
        RECT  8.685 6.255 9.135 6.705 ;
        RECT  2.205 6.255 2.655 6.705 ;
        END
    END rb
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER via ;
        RECT  6.525 4.725 6.795 4.995 ;
        RECT  3.915 4.725 4.185 4.995 ;
        LAYER metal2 ;
        RECT  6.435 4.635 6.885 5.085 ;
        RECT  3.825 4.680 6.885 5.040 ;
        RECT  3.825 4.635 4.275 5.085 ;
        LAYER metal1 ;
        RECT  6.435 4.635 6.885 5.085 ;
        RECT  3.825 4.635 4.275 5.085 ;
        END
    END ck
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 13.770 11.340 ;
        RECT  12.375 6.750 12.735 11.340 ;
        RECT  10.845 6.750 11.205 11.340 ;
        RECT  8.235 7.650 8.595 11.340 ;
        RECT  3.465 7.650 3.825 11.340 ;
        RECT  2.655 7.650 3.015 11.340 ;
        RECT  0.630 7.650 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 13.770 0.990 ;
        RECT  12.375 0.000 12.735 3.420 ;
        RECT  10.845 0.000 11.205 3.420 ;
        RECT  8.505 0.000 8.865 2.970 ;
        RECT  3.780 0.000 4.140 2.970 ;
        RECT  1.350 0.000 1.710 2.880 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  1.890 8.685 2.340 9.135 ;
        RECT  1.935 7.650 2.295 9.270 ;
        RECT  0.630 2.160 0.990 3.510 ;
        RECT  2.070 2.160 2.430 3.510 ;
        RECT  0.630 3.150 2.430 3.510 ;
        RECT  2.835 2.205 3.285 2.655 ;
        RECT  4.545 2.160 4.905 3.420 ;
        RECT  4.680 3.060 5.040 7.470 ;
        RECT  4.275 7.110 5.040 7.470 ;
        RECT  4.275 7.110 4.635 9.270 ;
        RECT  5.265 8.685 5.715 9.135 ;
        RECT  5.310 7.740 5.670 9.270 ;
        RECT  5.355 2.205 5.805 2.655 ;
        RECT  6.795 8.685 7.245 9.135 ;
        RECT  6.840 7.650 7.200 9.270 ;
        RECT  6.885 2.205 7.335 2.655 ;
        RECT  8.955 8.685 9.405 9.135 ;
        RECT  9.000 7.650 9.360 9.270 ;
        RECT  7.785 2.160 8.145 3.600 ;
        RECT  9.225 2.160 9.585 3.600 ;
        RECT  7.785 3.240 9.585 3.600 ;
        RECT  9.945 2.205 10.395 2.655 ;
        RECT  6.165 2.160 6.525 4.230 ;
        RECT  5.490 3.870 6.525 4.230 ;
        RECT  5.490 5.490 10.710 5.850 ;
        RECT  5.490 3.870 5.850 7.470 ;
        RECT  5.490 7.110 6.435 7.470 ;
        RECT  6.075 7.110 6.435 9.270 ;
        LAYER via ;
        RECT  1.980 8.775 2.250 9.045 ;
        RECT  2.925 2.295 3.195 2.565 ;
        RECT  5.355 8.775 5.625 9.045 ;
        RECT  5.445 2.295 5.715 2.565 ;
        RECT  6.885 8.775 7.155 9.045 ;
        RECT  6.975 2.295 7.245 2.565 ;
        RECT  9.045 8.775 9.315 9.045 ;
        RECT  10.035 2.295 10.305 2.565 ;
        LAYER metal2 ;
        RECT  1.890 8.730 5.715 9.090 ;
        RECT  1.890 8.685 2.340 9.135 ;
        RECT  5.265 8.685 5.715 9.135 ;
        RECT  2.835 2.250 5.805 2.610 ;
        RECT  2.835 2.205 3.285 2.655 ;
        RECT  5.355 2.205 5.805 2.655 ;
        RECT  6.795 8.730 9.405 9.090 ;
        RECT  6.795 8.685 7.245 9.135 ;
        RECT  8.955 8.685 9.405 9.135 ;
        RECT  6.885 2.250 10.395 2.610 ;
        RECT  6.885 2.205 7.335 2.655 ;
        RECT  9.945 2.205 10.395 2.655 ;
    END
END lrsp_4

MACRO lrsp_2
    CLASS CORE ;
    FOREIGN lrsp_2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.960 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER via ;
        RECT  6.525 4.725 6.795 4.995 ;
        RECT  3.915 4.725 4.185 4.995 ;
        LAYER metal2 ;
        RECT  6.435 4.635 6.885 5.085 ;
        RECT  3.825 4.680 6.885 5.040 ;
        RECT  3.825 4.635 4.275 5.085 ;
        LAYER metal1 ;
        RECT  6.435 4.635 6.885 5.085 ;
        RECT  3.825 4.635 4.275 5.085 ;
        END
    END ck
    PIN rb
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  8.775 6.345 9.045 6.615 ;
        RECT  2.295 6.345 2.565 6.615 ;
        LAYER metal2 ;
        RECT  8.685 6.255 9.135 6.705 ;
        RECT  2.205 6.300 9.135 6.660 ;
        RECT  2.205 6.255 2.655 6.705 ;
        LAYER metal1 ;
        RECT  8.685 6.255 9.135 6.705 ;
        RECT  2.205 6.255 2.655 6.705 ;
        END
    END rb
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.610 5.490 11.970 9.270 ;
        RECT  11.160 3.870 11.970 4.230 ;
        RECT  11.610 2.160 11.970 4.230 ;
        RECT  11.160 5.490 11.970 5.850 ;
        RECT  11.160 3.870 11.520 5.850 ;
        RECT  7.920 4.680 11.520 5.040 ;
        END
    END q
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip
    PIN s
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  7.155 3.915 7.425 4.185 ;
        RECT  1.485 3.915 1.755 4.185 ;
        LAYER metal2 ;
        RECT  7.065 3.825 7.515 4.275 ;
        RECT  1.395 3.870 7.515 4.230 ;
        RECT  1.395 3.825 1.845 4.275 ;
        LAYER metal1 ;
        RECT  7.065 3.825 7.515 4.275 ;
        RECT  1.395 3.825 1.845 4.275 ;
        END
    END s
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 12.960 11.340 ;
        RECT  10.845 6.750 11.205 11.340 ;
        RECT  8.235 7.650 8.595 11.340 ;
        RECT  3.465 7.650 3.825 11.340 ;
        RECT  2.655 7.650 3.015 11.340 ;
        RECT  0.630 7.650 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 12.960 0.990 ;
        RECT  10.845 0.000 11.205 3.420 ;
        RECT  8.505 0.000 8.865 2.970 ;
        RECT  3.780 0.000 4.140 2.970 ;
        RECT  1.350 0.000 1.710 2.880 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  1.890 8.685 2.340 9.135 ;
        RECT  1.935 7.650 2.295 9.270 ;
        RECT  0.630 2.160 0.990 3.510 ;
        RECT  2.070 2.160 2.430 3.510 ;
        RECT  0.630 3.150 2.430 3.510 ;
        RECT  2.835 2.205 3.285 2.655 ;
        RECT  4.545 2.160 4.905 3.420 ;
        RECT  4.680 3.060 5.040 7.470 ;
        RECT  4.275 7.110 5.040 7.470 ;
        RECT  4.275 7.110 4.635 9.270 ;
        RECT  5.265 8.685 5.715 9.135 ;
        RECT  5.310 7.740 5.670 9.270 ;
        RECT  5.355 2.205 5.805 2.655 ;
        RECT  6.795 8.685 7.245 9.135 ;
        RECT  6.840 7.650 7.200 9.270 ;
        RECT  6.885 2.205 7.335 2.655 ;
        RECT  8.955 8.685 9.405 9.135 ;
        RECT  9.000 7.650 9.360 9.270 ;
        RECT  7.785 2.160 8.145 3.600 ;
        RECT  9.225 2.160 9.585 3.600 ;
        RECT  7.785 3.240 9.585 3.600 ;
        RECT  9.945 2.205 10.395 2.655 ;
        RECT  6.165 2.160 6.525 4.230 ;
        RECT  5.490 3.870 6.525 4.230 ;
        RECT  5.490 5.490 10.710 5.850 ;
        RECT  5.490 3.870 5.850 7.470 ;
        RECT  5.490 7.110 6.435 7.470 ;
        RECT  6.075 7.110 6.435 9.270 ;
        LAYER via ;
        RECT  1.980 8.775 2.250 9.045 ;
        RECT  2.925 2.295 3.195 2.565 ;
        RECT  5.355 8.775 5.625 9.045 ;
        RECT  5.445 2.295 5.715 2.565 ;
        RECT  6.885 8.775 7.155 9.045 ;
        RECT  6.975 2.295 7.245 2.565 ;
        RECT  9.045 8.775 9.315 9.045 ;
        RECT  10.035 2.295 10.305 2.565 ;
        LAYER metal2 ;
        RECT  1.890 8.730 5.715 9.090 ;
        RECT  1.890 8.685 2.340 9.135 ;
        RECT  5.265 8.685 5.715 9.135 ;
        RECT  2.835 2.250 5.805 2.610 ;
        RECT  2.835 2.205 3.285 2.655 ;
        RECT  5.355 2.205 5.805 2.655 ;
        RECT  6.795 8.730 9.405 9.090 ;
        RECT  6.795 8.685 7.245 9.135 ;
        RECT  8.955 8.685 9.405 9.135 ;
        RECT  6.885 2.250 10.395 2.610 ;
        RECT  6.885 2.205 7.335 2.655 ;
        RECT  9.945 2.205 10.395 2.655 ;
    END
END lrsp_2

MACRO lrsp_1
    CLASS CORE ;
    FOREIGN lrsp_1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.960 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER via ;
        RECT  6.525 4.725 6.795 4.995 ;
        RECT  3.915 4.725 4.185 4.995 ;
        LAYER metal2 ;
        RECT  6.435 4.635 6.885 5.085 ;
        RECT  3.825 4.680 6.885 5.040 ;
        RECT  3.825 4.635 4.275 5.085 ;
        LAYER metal1 ;
        RECT  6.435 4.635 6.885 5.085 ;
        RECT  3.825 4.635 4.275 5.085 ;
        END
    END ck
    PIN rb
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  8.775 6.345 9.045 6.615 ;
        RECT  2.295 6.345 2.565 6.615 ;
        LAYER metal2 ;
        RECT  8.685 6.255 9.135 6.705 ;
        RECT  2.205 6.300 9.135 6.660 ;
        RECT  2.205 6.255 2.655 6.705 ;
        LAYER metal1 ;
        RECT  8.685 6.255 9.135 6.705 ;
        RECT  2.205 6.255 2.655 6.705 ;
        END
    END rb
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.610 5.490 11.970 9.270 ;
        RECT  11.160 3.870 11.970 4.230 ;
        RECT  11.610 2.160 11.970 4.230 ;
        RECT  11.160 5.490 11.970 5.850 ;
        RECT  11.160 3.870 11.520 5.850 ;
        RECT  7.920 4.680 11.520 5.040 ;
        END
    END q
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip
    PIN s
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  7.155 3.915 7.425 4.185 ;
        RECT  1.485 3.915 1.755 4.185 ;
        LAYER metal2 ;
        RECT  7.065 3.825 7.515 4.275 ;
        RECT  1.395 3.870 7.515 4.230 ;
        RECT  1.395 3.825 1.845 4.275 ;
        LAYER metal1 ;
        RECT  7.065 3.825 7.515 4.275 ;
        RECT  1.395 3.825 1.845 4.275 ;
        END
    END s
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 12.960 0.990 ;
        RECT  10.845 0.000 11.205 2.970 ;
        RECT  8.505 0.000 8.865 2.970 ;
        RECT  3.780 0.000 4.140 2.970 ;
        RECT  1.350 0.000 1.710 2.880 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 12.960 11.340 ;
        RECT  10.845 7.650 11.205 11.340 ;
        RECT  8.235 7.650 8.595 11.340 ;
        RECT  3.465 7.650 3.825 11.340 ;
        RECT  2.655 7.650 3.015 11.340 ;
        RECT  0.630 7.650 0.990 11.340 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  1.890 8.685 2.340 9.135 ;
        RECT  1.935 7.650 2.295 9.270 ;
        RECT  0.630 2.160 0.990 3.510 ;
        RECT  2.070 2.160 2.430 3.510 ;
        RECT  0.630 3.150 2.430 3.510 ;
        RECT  2.835 2.205 3.285 2.655 ;
        RECT  4.545 2.160 4.905 3.420 ;
        RECT  4.680 3.060 5.040 7.470 ;
        RECT  4.275 7.110 5.040 7.470 ;
        RECT  4.275 7.110 4.635 9.270 ;
        RECT  5.265 8.685 5.715 9.135 ;
        RECT  5.310 7.740 5.670 9.270 ;
        RECT  5.355 2.205 5.805 2.655 ;
        RECT  6.795 8.685 7.245 9.135 ;
        RECT  6.840 7.650 7.200 9.270 ;
        RECT  6.885 2.205 7.335 2.655 ;
        RECT  8.955 8.685 9.405 9.135 ;
        RECT  9.000 7.650 9.360 9.270 ;
        RECT  7.785 2.160 8.145 3.600 ;
        RECT  9.225 2.160 9.585 3.600 ;
        RECT  7.785 3.240 9.585 3.600 ;
        RECT  9.945 2.205 10.395 2.655 ;
        RECT  6.165 2.160 6.525 4.230 ;
        RECT  5.490 3.870 6.525 4.230 ;
        RECT  5.490 5.490 10.710 5.850 ;
        RECT  5.490 3.870 5.850 7.470 ;
        RECT  5.490 7.110 6.435 7.470 ;
        RECT  6.075 7.110 6.435 9.270 ;
        LAYER via ;
        RECT  1.980 8.775 2.250 9.045 ;
        RECT  2.925 2.295 3.195 2.565 ;
        RECT  5.355 8.775 5.625 9.045 ;
        RECT  5.445 2.295 5.715 2.565 ;
        RECT  6.885 8.775 7.155 9.045 ;
        RECT  6.975 2.295 7.245 2.565 ;
        RECT  9.045 8.775 9.315 9.045 ;
        RECT  10.035 2.295 10.305 2.565 ;
        LAYER metal2 ;
        RECT  1.890 8.730 5.715 9.090 ;
        RECT  1.890 8.685 2.340 9.135 ;
        RECT  5.265 8.685 5.715 9.135 ;
        RECT  2.835 2.250 5.805 2.610 ;
        RECT  2.835 2.205 3.285 2.655 ;
        RECT  5.355 2.205 5.805 2.655 ;
        RECT  6.795 8.730 9.405 9.090 ;
        RECT  6.795 8.685 7.245 9.135 ;
        RECT  8.955 8.685 9.405 9.135 ;
        RECT  6.885 2.250 10.395 2.610 ;
        RECT  6.885 2.205 7.335 2.655 ;
        RECT  9.945 2.205 10.395 2.655 ;
    END
END lrsp_1

MACRO lrp_4
    CLASS CORE ;
    FOREIGN lrp_4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.150 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 4.680 0.990 5.040 ;
        END
    END ip
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER via ;
        RECT  5.940 4.725 6.210 4.995 ;
        RECT  3.105 4.725 3.375 4.995 ;
        LAYER metal2 ;
        RECT  5.850 4.635 6.300 5.085 ;
        RECT  3.015 4.680 6.300 5.040 ;
        RECT  3.015 4.635 3.465 5.085 ;
        LAYER metal1 ;
        RECT  5.850 4.635 6.300 5.085 ;
        RECT  3.015 4.635 3.465 5.085 ;
        RECT  3.060 4.635 3.420 5.850 ;
        END
    END ck
    PIN rb
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  7.965 6.345 8.235 6.615 ;
        RECT  2.295 6.345 2.565 6.615 ;
        LAYER metal2 ;
        RECT  7.875 6.255 8.325 6.705 ;
        RECT  2.205 6.300 8.325 6.660 ;
        RECT  2.205 6.255 2.655 6.705 ;
        LAYER metal1 ;
        RECT  7.875 6.255 8.325 6.705 ;
        RECT  2.205 6.255 2.655 6.705 ;
        END
    END rb
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.350 3.870 10.710 5.850 ;
        RECT  10.080 5.490 10.440 9.270 ;
        RECT  7.110 4.680 10.710 5.040 ;
        RECT  10.080 2.160 10.440 4.230 ;
        END
    END q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 12.150 11.340 ;
        RECT  10.845 6.750 11.205 11.340 ;
        RECT  9.315 6.750 9.675 11.340 ;
        RECT  7.020 7.740 7.380 11.340 ;
        RECT  2.925 7.650 3.285 11.340 ;
        RECT  2.115 7.650 2.475 11.340 ;
        RECT  0.630 7.650 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 12.150 0.990 ;
        RECT  10.845 0.000 11.205 3.420 ;
        RECT  9.315 0.000 9.675 3.420 ;
        RECT  6.885 0.000 7.245 2.970 ;
        RECT  2.835 0.000 3.195 2.970 ;
        RECT  0.630 0.000 0.990 2.970 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  1.305 8.685 1.755 9.135 ;
        RECT  1.350 7.650 1.710 9.270 ;
        RECT  1.890 2.205 2.340 2.655 ;
        RECT  3.600 2.160 3.960 3.420 ;
        RECT  3.870 3.060 4.230 6.660 ;
        RECT  3.690 6.300 4.050 9.270 ;
        RECT  4.410 2.205 4.860 2.655 ;
        RECT  4.680 8.685 5.130 9.135 ;
        RECT  4.725 7.650 5.085 9.270 ;
        RECT  6.255 7.110 8.190 7.470 ;
        RECT  6.255 7.110 6.615 9.270 ;
        RECT  7.830 7.110 8.190 9.270 ;
        RECT  5.985 2.160 6.345 3.825 ;
        RECT  8.325 2.160 8.685 3.825 ;
        RECT  5.985 3.465 8.685 3.825 ;
        RECT  5.220 2.160 5.580 4.230 ;
        RECT  4.680 3.870 5.580 4.230 ;
        RECT  4.680 5.490 9.495 5.850 ;
        RECT  4.680 3.870 5.040 6.660 ;
        RECT  4.680 6.300 5.850 6.660 ;
        RECT  5.490 6.300 5.850 9.270 ;
        LAYER via ;
        RECT  1.395 8.775 1.665 9.045 ;
        RECT  1.980 2.295 2.250 2.565 ;
        RECT  4.500 2.295 4.770 2.565 ;
        RECT  4.770 8.775 5.040 9.045 ;
        LAYER metal2 ;
        RECT  1.890 2.250 4.860 2.610 ;
        RECT  1.890 2.205 2.340 2.655 ;
        RECT  4.410 2.205 4.860 2.655 ;
        RECT  1.305 8.730 5.130 9.090 ;
        RECT  1.305 8.685 1.755 9.135 ;
        RECT  4.680 8.685 5.130 9.135 ;
    END
END lrp_4

MACRO lrp_2
    CLASS CORE ;
    FOREIGN lrp_2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.340 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.350 3.870 10.710 5.850 ;
        RECT  10.080 5.490 10.440 9.270 ;
        RECT  7.110 4.680 10.710 5.040 ;
        RECT  10.080 2.160 10.440 4.230 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  7.965 6.345 8.235 6.615 ;
        RECT  2.295 6.345 2.565 6.615 ;
        LAYER metal2 ;
        RECT  7.875 6.255 8.325 6.705 ;
        RECT  2.205 6.300 8.325 6.660 ;
        RECT  2.205 6.255 2.655 6.705 ;
        LAYER metal1 ;
        RECT  7.875 6.255 8.325 6.705 ;
        RECT  2.205 6.255 2.655 6.705 ;
        END
    END rb
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER via ;
        RECT  5.940 4.725 6.210 4.995 ;
        RECT  3.105 4.725 3.375 4.995 ;
        LAYER metal2 ;
        RECT  5.850 4.635 6.300 5.085 ;
        RECT  3.015 4.680 6.300 5.040 ;
        RECT  3.015 4.635 3.465 5.085 ;
        LAYER metal1 ;
        RECT  5.850 4.635 6.300 5.085 ;
        RECT  3.015 4.635 3.465 5.085 ;
        RECT  3.060 4.635 3.420 5.850 ;
        END
    END ck
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 4.680 0.990 5.040 ;
        END
    END ip
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 11.340 11.340 ;
        RECT  9.315 6.750 9.675 11.340 ;
        RECT  7.020 7.740 7.380 11.340 ;
        RECT  2.925 7.650 3.285 11.340 ;
        RECT  2.115 7.650 2.475 11.340 ;
        RECT  0.630 7.650 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 11.340 0.990 ;
        RECT  9.315 0.000 9.675 3.420 ;
        RECT  6.885 0.000 7.245 2.970 ;
        RECT  2.835 0.000 3.195 2.970 ;
        RECT  0.630 0.000 0.990 2.970 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  1.305 8.685 1.755 9.135 ;
        RECT  1.350 7.650 1.710 9.270 ;
        RECT  1.890 2.205 2.340 2.655 ;
        RECT  3.600 2.160 3.960 3.420 ;
        RECT  3.870 3.060 4.230 6.660 ;
        RECT  3.690 6.300 4.050 9.270 ;
        RECT  4.410 2.205 4.860 2.655 ;
        RECT  4.680 8.685 5.130 9.135 ;
        RECT  4.725 7.650 5.085 9.270 ;
        RECT  6.255 7.110 8.190 7.470 ;
        RECT  6.255 7.110 6.615 9.270 ;
        RECT  7.830 7.110 8.190 9.270 ;
        RECT  5.985 2.160 6.345 3.825 ;
        RECT  8.325 2.160 8.685 3.825 ;
        RECT  5.985 3.465 8.685 3.825 ;
        RECT  5.220 2.160 5.580 4.230 ;
        RECT  4.680 3.870 5.580 4.230 ;
        RECT  4.680 5.490 9.495 5.850 ;
        RECT  4.680 3.870 5.040 6.660 ;
        RECT  4.680 6.300 5.850 6.660 ;
        RECT  5.490 6.300 5.850 9.270 ;
        LAYER via ;
        RECT  1.395 8.775 1.665 9.045 ;
        RECT  1.980 2.295 2.250 2.565 ;
        RECT  4.500 2.295 4.770 2.565 ;
        RECT  4.770 8.775 5.040 9.045 ;
        LAYER metal2 ;
        RECT  1.890 2.250 4.860 2.610 ;
        RECT  1.890 2.205 2.340 2.655 ;
        RECT  4.410 2.205 4.860 2.655 ;
        RECT  1.305 8.730 5.130 9.090 ;
        RECT  1.305 8.685 1.755 9.135 ;
        RECT  4.680 8.685 5.130 9.135 ;
    END
END lrp_2

MACRO lrp_1
    CLASS CORE ;
    FOREIGN lrp_1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.340 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.350 3.060 10.710 7.470 ;
        RECT  10.080 7.110 10.440 9.270 ;
        RECT  7.110 4.680 10.710 5.040 ;
        RECT  10.080 2.160 10.440 3.420 ;
        END
    END q
    PIN rb
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  7.965 6.345 8.235 6.615 ;
        RECT  2.295 6.345 2.565 6.615 ;
        LAYER metal2 ;
        RECT  7.875 6.255 8.325 6.705 ;
        RECT  2.205 6.300 8.325 6.660 ;
        RECT  2.205 6.255 2.655 6.705 ;
        LAYER metal1 ;
        RECT  7.875 6.255 8.325 6.705 ;
        RECT  2.205 6.255 2.655 6.705 ;
        END
    END rb
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER via ;
        RECT  5.940 4.725 6.210 4.995 ;
        RECT  3.105 4.725 3.375 4.995 ;
        LAYER metal2 ;
        RECT  5.850 4.635 6.300 5.085 ;
        RECT  3.015 4.680 6.300 5.040 ;
        RECT  3.015 4.635 3.465 5.085 ;
        LAYER metal1 ;
        RECT  5.850 4.635 6.300 5.085 ;
        RECT  3.015 4.635 3.465 5.085 ;
        RECT  3.060 4.635 3.420 5.850 ;
        END
    END ck
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 4.680 0.990 5.040 ;
        END
    END ip
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 11.340 0.990 ;
        RECT  9.315 0.000 9.675 2.970 ;
        RECT  6.885 0.000 7.245 2.970 ;
        RECT  2.835 0.000 3.195 2.970 ;
        RECT  0.630 0.000 0.990 2.970 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 11.340 11.340 ;
        RECT  9.315 7.650 9.675 11.340 ;
        RECT  7.020 7.740 7.380 11.340 ;
        RECT  2.925 7.650 3.285 11.340 ;
        RECT  2.115 7.650 2.475 11.340 ;
        RECT  0.630 7.650 0.990 11.340 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  1.305 8.685 1.755 9.135 ;
        RECT  1.350 7.650 1.710 9.270 ;
        RECT  1.890 2.205 2.340 2.655 ;
        RECT  3.600 2.160 3.960 3.420 ;
        RECT  3.870 3.060 4.230 6.660 ;
        RECT  3.690 6.300 4.050 9.270 ;
        RECT  4.410 2.205 4.860 2.655 ;
        RECT  4.680 8.685 5.130 9.135 ;
        RECT  4.725 7.650 5.085 9.270 ;
        RECT  6.255 7.110 8.190 7.470 ;
        RECT  6.255 7.110 6.615 9.270 ;
        RECT  7.830 7.110 8.190 9.270 ;
        RECT  5.985 2.160 6.345 3.825 ;
        RECT  8.325 2.160 8.685 3.825 ;
        RECT  5.985 3.465 8.685 3.825 ;
        RECT  5.220 2.160 5.580 4.230 ;
        RECT  4.680 3.870 5.580 4.230 ;
        RECT  4.680 5.490 9.495 5.850 ;
        RECT  4.680 3.870 5.040 6.660 ;
        RECT  4.680 6.300 5.850 6.660 ;
        RECT  5.490 6.300 5.850 9.270 ;
        LAYER via ;
        RECT  1.395 8.775 1.665 9.045 ;
        RECT  1.980 2.295 2.250 2.565 ;
        RECT  4.500 2.295 4.770 2.565 ;
        RECT  4.770 8.775 5.040 9.045 ;
        LAYER metal2 ;
        RECT  1.890 2.250 4.860 2.610 ;
        RECT  1.890 2.205 2.340 2.655 ;
        RECT  4.410 2.205 4.860 2.655 ;
        RECT  1.305 8.730 5.130 9.090 ;
        RECT  1.305 8.685 1.755 9.135 ;
        RECT  4.680 8.685 5.130 9.135 ;
    END
END lrp_1

MACRO lp_2
    CLASS CORE ;
    FOREIGN lp_2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.100 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER metal1 ;
        RECT  1.440 3.870 3.420 4.230 ;
        END
    END ck
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 4.680 2.610 5.040 ;
        END
    END ip
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.670 6.300 6.660 6.660 ;
        RECT  6.300 3.870 6.660 6.660 ;
        RECT  4.680 3.870 6.660 4.230 ;
        RECT  5.670 6.300 6.030 9.270 ;
        RECT  5.670 2.160 6.030 4.230 ;
        END
    END q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 8.100 11.340 ;
        RECT  6.480 6.975 6.840 11.340 ;
        RECT  4.905 6.975 5.265 11.340 ;
        RECT  2.025 6.975 2.385 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 8.100 0.990 ;
        RECT  6.525 0.000 6.885 3.420 ;
        RECT  4.860 0.000 5.220 3.420 ;
        RECT  2.025 0.000 2.385 3.420 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  1.215 2.160 1.575 3.420 ;
        RECT  0.630 3.060 1.575 3.420 ;
        RECT  0.630 3.060 0.990 6.660 ;
        RECT  0.630 6.300 3.420 6.660 ;
        RECT  1.215 6.300 1.575 9.270 ;
        RECT  1.440 5.490 4.230 5.850 ;
        RECT  3.375 2.160 3.735 3.600 ;
        RECT  3.375 3.240 4.230 3.600 ;
        RECT  3.870 3.240 4.230 5.040 ;
        RECT  3.870 4.680 5.850 5.040 ;
        RECT  4.860 4.680 5.220 6.660 ;
        RECT  4.230 6.300 5.220 6.660 ;
        RECT  4.230 6.300 4.590 7.290 ;
        RECT  3.465 6.930 4.590 7.290 ;
        RECT  3.465 6.930 3.825 9.270 ;
    END
END lp_2

MACRO lp_1
    CLASS CORE ;
    FOREIGN lp_1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.290 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.445 6.300 6.660 6.660 ;
        RECT  6.300 3.870 6.660 6.660 ;
        RECT  4.680 3.870 6.660 4.230 ;
        RECT  5.445 6.300 5.805 9.270 ;
        RECT  5.445 2.160 5.805 4.230 ;
        END
    END q
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 4.680 2.610 5.040 ;
        END
    END ip
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER metal1 ;
        RECT  1.440 3.870 3.195 4.230 ;
        END
    END ck
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 7.290 0.990 ;
        RECT  6.300 0.000 6.660 2.790 ;
        RECT  4.635 0.000 4.995 2.790 ;
        RECT  1.800 0.000 2.160 2.790 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 7.290 11.340 ;
        RECT  6.255 8.010 6.615 11.340 ;
        RECT  4.680 8.010 5.040 11.340 ;
        RECT  1.800 8.010 2.160 11.340 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  0.990 2.160 1.350 3.420 ;
        RECT  0.630 3.060 0.990 7.470 ;
        RECT  0.630 7.110 3.195 7.470 ;
        RECT  0.990 7.110 1.350 9.270 ;
        RECT  1.440 5.490 4.005 5.850 ;
        RECT  3.150 2.160 3.510 3.600 ;
        RECT  3.150 3.240 4.005 3.600 ;
        RECT  3.645 3.240 4.005 5.040 ;
        RECT  3.645 4.680 5.625 5.040 ;
        RECT  4.635 4.680 4.995 6.660 ;
        RECT  4.005 6.300 4.995 6.660 ;
        RECT  4.005 6.300 4.365 8.190 ;
        RECT  3.240 7.830 4.365 8.190 ;
        RECT  3.240 7.830 3.600 9.270 ;
    END
END lp_1

MACRO jkrp_2
    CLASS CORE ;
    FOREIGN jkrp_2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 27.540 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN j
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END j
    PIN k
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  3.870 6.300 4.230 6.660 ;
        END
    END k
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER metal1 ;
        RECT  7.920 4.680 8.280 5.040 ;
        END
    END ck
    PIN rb
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  20.340 5.535 20.610 5.805 ;
        RECT  16.065 5.535 16.335 5.805 ;
        LAYER metal2 ;
        RECT  20.250 5.445 20.700 5.895 ;
        RECT  15.975 5.490 20.700 5.850 ;
        RECT  15.975 5.445 16.425 5.895 ;
        LAYER metal1 ;
        RECT  20.250 5.445 20.700 5.895 ;
        RECT  15.975 5.445 16.425 5.895 ;
        END
    END rb
    PIN qb
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  24.795 4.500 25.290 6.300 ;
        RECT  24.795 2.160 25.155 9.270 ;
        END
    END qb
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  26.280 4.275 26.910 6.075 ;
        RECT  26.280 2.160 26.640 9.270 ;
        END
    END q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 27.540 11.340 ;
        RECT  25.515 6.750 25.875 11.340 ;
        RECT  24.030 6.750 24.390 11.340 ;
        RECT  22.545 8.010 22.905 11.340 ;
        RECT  21.825 8.010 22.185 11.340 ;
        RECT  20.295 8.010 20.655 11.340 ;
        RECT  16.020 8.010 16.380 11.340 ;
        RECT  14.490 8.010 14.850 11.340 ;
        RECT  12.735 8.010 13.095 11.340 ;
        RECT  9.225 8.010 9.585 11.340 ;
        RECT  7.740 8.010 8.100 11.340 ;
        RECT  3.015 8.010 3.375 11.340 ;
        RECT  0.630 8.010 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 27.540 0.990 ;
        RECT  25.515 0.000 25.875 3.420 ;
        RECT  24.030 0.000 24.390 3.420 ;
        RECT  22.545 0.000 22.905 2.655 ;
        RECT  20.295 0.000 20.655 2.655 ;
        RECT  14.490 0.000 14.850 2.655 ;
        RECT  12.735 0.000 13.095 2.655 ;
        RECT  9.225 0.000 9.585 2.655 ;
        RECT  7.740 0.000 8.100 2.655 ;
        RECT  5.265 0.000 5.625 2.655 ;
        RECT  2.205 0.000 2.565 2.790 ;
        RECT  0.630 0.000 0.990 2.790 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  2.205 8.685 2.655 9.135 ;
        RECT  2.205 8.010 2.565 9.270 ;
        RECT  2.205 3.825 2.655 4.275 ;
        RECT  1.395 5.490 3.780 5.850 ;
        RECT  1.395 2.295 1.755 9.270 ;
        RECT  3.690 8.685 4.140 9.135 ;
        RECT  3.735 8.010 4.095 9.270 ;
        RECT  5.220 8.685 5.670 9.135 ;
        RECT  5.265 8.010 5.625 9.270 ;
        RECT  5.220 3.015 5.670 3.465 ;
        RECT  3.735 2.250 4.095 5.040 ;
        RECT  3.735 4.680 6.435 5.040 ;
        RECT  4.545 7.110 6.435 7.470 ;
        RECT  4.545 7.110 4.905 9.270 ;
        RECT  6.075 2.160 6.435 9.270 ;
        RECT  6.795 5.445 7.245 5.895 ;
        RECT  6.840 2.160 7.200 9.270 ;
        RECT  7.470 7.065 7.920 7.515 ;
        RECT  7.470 3.555 8.865 3.915 ;
        RECT  8.505 2.160 8.865 4.365 ;
        RECT  8.730 4.005 9.090 5.850 ;
        RECT  8.505 5.490 9.720 5.850 ;
        RECT  8.505 6.255 8.955 6.705 ;
        RECT  8.505 5.490 8.865 9.270 ;
        RECT  9.990 2.160 10.350 3.420 ;
        RECT  10.350 3.060 10.710 4.230 ;
        RECT  9.945 4.635 10.395 5.085 ;
        RECT  9.945 7.065 10.395 7.515 ;
        RECT  9.990 3.870 10.350 9.270 ;
        RECT  10.935 5.445 11.385 5.895 ;
        RECT  10.980 2.160 11.340 9.270 ;
        RECT  12.465 6.255 12.915 6.705 ;
        RECT  11.745 7.110 13.860 7.470 ;
        RECT  11.745 2.160 12.105 9.270 ;
        RECT  13.500 2.160 13.860 9.270 ;
        RECT  14.355 5.445 14.805 5.895 ;
        RECT  16.245 6.255 16.695 6.705 ;
        RECT  16.245 4.635 16.695 5.085 ;
        RECT  16.020 2.160 16.380 4.230 ;
        RECT  15.255 3.870 17.370 4.230 ;
        RECT  14.220 6.300 15.615 6.660 ;
        RECT  15.255 3.870 15.615 9.270 ;
        RECT  17.010 2.160 17.370 9.270 ;
        RECT  17.730 4.635 18.180 5.085 ;
        RECT  17.775 5.490 18.900 5.850 ;
        RECT  17.775 2.160 18.135 9.270 ;
        RECT  18.540 2.160 18.900 9.270 ;
        RECT  20.025 7.065 20.475 7.515 ;
        RECT  21.825 2.160 22.185 4.230 ;
        RECT  21.060 3.870 22.185 4.230 ;
        RECT  21.060 3.825 21.510 4.275 ;
        RECT  19.305 6.300 21.465 6.660 ;
        RECT  19.305 2.160 19.665 9.270 ;
        RECT  21.105 3.825 21.465 9.270 ;
        RECT  22.455 4.635 22.905 5.085 ;
        RECT  23.265 3.015 23.715 3.465 ;
        RECT  23.310 5.490 24.390 5.850 ;
        RECT  21.870 7.110 23.670 7.470 ;
        RECT  23.310 2.160 23.670 9.270 ;
        RECT  25.470 3.825 25.920 4.275 ;
        LAYER via ;
        RECT  2.295 8.775 2.565 9.045 ;
        RECT  2.295 3.915 2.565 4.185 ;
        RECT  3.780 8.775 4.050 9.045 ;
        RECT  5.310 8.775 5.580 9.045 ;
        RECT  5.310 3.105 5.580 3.375 ;
        RECT  6.885 5.535 7.155 5.805 ;
        RECT  7.560 7.155 7.830 7.425 ;
        RECT  8.595 6.345 8.865 6.615 ;
        RECT  10.035 7.155 10.305 7.425 ;
        RECT  10.035 4.725 10.305 4.995 ;
        RECT  11.025 5.535 11.295 5.805 ;
        RECT  12.555 6.345 12.825 6.615 ;
        RECT  14.445 5.535 14.715 5.805 ;
        RECT  16.335 6.345 16.605 6.615 ;
        RECT  16.335 4.725 16.605 4.995 ;
        RECT  17.820 4.725 18.090 4.995 ;
        RECT  20.115 7.155 20.385 7.425 ;
        RECT  21.150 3.915 21.420 4.185 ;
        RECT  22.545 4.725 22.815 4.995 ;
        RECT  23.355 3.105 23.625 3.375 ;
        RECT  25.560 3.915 25.830 4.185 ;
        LAYER metal2 ;
        RECT  2.205 8.730 5.670 9.090 ;
        RECT  2.205 8.685 2.655 9.135 ;
        RECT  3.690 8.685 4.140 9.135 ;
        RECT  5.220 8.685 5.670 9.135 ;
        RECT  6.795 5.490 14.805 5.850 ;
        RECT  6.795 5.445 7.245 5.895 ;
        RECT  10.935 5.445 11.385 5.895 ;
        RECT  14.355 5.445 14.805 5.895 ;
        RECT  8.505 6.300 16.695 6.660 ;
        RECT  8.505 6.255 8.955 6.705 ;
        RECT  12.465 6.255 12.915 6.705 ;
        RECT  16.245 6.255 16.695 6.705 ;
        RECT  9.945 4.680 16.695 5.040 ;
        RECT  9.945 4.635 10.395 5.085 ;
        RECT  16.245 4.635 16.695 5.085 ;
        RECT  7.470 7.110 20.475 7.470 ;
        RECT  7.470 7.065 7.920 7.515 ;
        RECT  9.945 7.065 10.395 7.515 ;
        RECT  20.025 7.065 20.475 7.515 ;
        RECT  17.730 4.680 22.905 5.040 ;
        RECT  17.730 4.635 18.180 5.085 ;
        RECT  22.455 4.635 22.905 5.085 ;
        RECT  5.220 3.060 23.715 3.420 ;
        RECT  5.220 3.015 5.670 3.465 ;
        RECT  23.265 3.015 23.715 3.465 ;
        RECT  2.205 3.870 25.920 4.230 ;
        RECT  2.205 3.825 2.655 4.275 ;
        RECT  21.060 3.825 21.510 4.275 ;
        RECT  25.470 3.825 25.920 4.275 ;
    END
END jkrp_2

MACRO invzp_4
    CLASS CORE ;
    FOREIGN invzp_4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN c
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 5.490 3.420 5.850 ;
        RECT  1.440 4.680 1.800 5.850 ;
        END
    END c
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  3.060 4.680 3.420 5.040 ;
        END
    END ip
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.970 6.120 4.230 6.480 ;
        RECT  3.870 3.555 4.230 6.480 ;
        RECT  3.555 3.105 3.915 3.915 ;
        RECT  2.880 3.105 3.915 3.465 ;
        RECT  2.970 6.120 3.330 9.270 ;
        RECT  2.880 2.160 3.240 3.465 ;
        END
    END op
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 5.670 11.340 ;
        RECT  4.320 6.750 4.680 11.340 ;
        RECT  1.620 6.750 1.980 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 5.670 0.990 ;
        RECT  4.230 0.000 4.590 3.240 ;
        RECT  1.530 0.000 1.890 3.420 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  0.630 3.870 3.195 4.230 ;
        RECT  0.630 2.160 0.990 9.270 ;
    END
END invzp_4

MACRO invzp_2
    CLASS CORE ;
    FOREIGN invzp_2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.860 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.970 6.120 4.230 6.480 ;
        RECT  3.870 3.105 4.230 6.480 ;
        RECT  2.880 3.105 4.230 3.465 ;
        RECT  2.970 6.120 3.330 9.270 ;
        RECT  2.880 2.160 3.240 3.465 ;
        END
    END op
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 4.680 2.610 5.040 ;
        END
    END ip
    PIN c
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 5.490 3.420 5.850 ;
        END
    END c
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 4.860 0.990 ;
        RECT  1.530 0.000 1.890 3.420 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 4.860 11.340 ;
        RECT  1.620 6.750 1.980 11.340 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  0.630 3.870 3.195 4.230 ;
        RECT  0.630 2.160 0.990 9.270 ;
    END
END invzp_2

MACRO invzp_1
    CLASS CORE ;
    FOREIGN invzp_1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.050 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.060 3.105 3.420 8.235 ;
        RECT  2.970 7.875 3.330 9.270 ;
        RECT  2.880 2.160 3.240 3.465 ;
        END
    END op
    PIN c
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 5.490 2.610 7.470 ;
        RECT  1.440 5.490 2.610 5.850 ;
        END
    END c
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 4.680 2.610 5.040 ;
        END
    END ip
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 4.050 0.990 ;
        RECT  1.530 0.000 1.890 2.790 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 4.050 11.340 ;
        RECT  1.620 8.010 1.980 11.340 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  0.630 3.870 2.610 4.230 ;
        RECT  0.630 2.160 0.990 9.270 ;
    END
END invzp_1

MACRO inv_4
    CLASS CORE ;
    FOREIGN inv_4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.240 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.395 5.490 2.610 5.850 ;
        RECT  2.250 3.870 2.610 5.850 ;
        RECT  1.395 3.870 2.610 4.230 ;
        RECT  1.395 5.490 1.755 9.270 ;
        RECT  1.395 2.160 1.755 4.230 ;
        END
    END op
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 4.680 0.990 5.040 ;
        END
    END ip
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 3.240 11.340 ;
        RECT  2.115 6.750 2.475 11.340 ;
        RECT  0.630 6.750 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 3.240 0.990 ;
        RECT  2.115 0.000 2.475 3.420 ;
        RECT  0.630 0.000 0.990 3.420 ;
        END
    END gnd!
END inv_4

MACRO inv_2
    CLASS CORE ;
    FOREIGN inv_2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.430 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 4.680 0.990 5.040 ;
        END
    END ip
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.440 3.285 1.800 6.660 ;
        RECT  1.395 6.300 1.755 9.270 ;
        RECT  1.395 2.160 1.755 3.645 ;
        END
    END op
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 2.430 0.990 ;
        RECT  0.630 0.000 0.990 3.420 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 2.430 11.340 ;
        RECT  0.630 6.750 0.990 11.340 ;
        END
    END vdd!
END inv_2

MACRO inv_1
    CLASS CORE ;
    FOREIGN inv_1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.430 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 4.680 0.990 5.040 ;
        END
    END ip
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.440 3.060 1.800 6.660 ;
        RECT  1.395 6.300 1.755 9.270 ;
        RECT  1.395 2.160 1.755 3.420 ;
        END
    END op
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 2.430 0.990 ;
        RECT  0.630 0.000 0.990 2.790 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 2.430 11.340 ;
        RECT  0.630 8.010 0.990 11.340 ;
        END
    END vdd!
END inv_1

MACRO fulladder
    CLASS CORE ;
    FOREIGN fulladder 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.820 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN a
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  12.960 6.345 13.230 6.615 ;
        RECT  8.640 6.345 8.910 6.615 ;
        RECT  4.410 6.345 4.680 6.615 ;
        RECT  1.485 6.345 1.755 6.615 ;
        LAYER metal2 ;
        RECT  12.870 6.255 13.320 6.705 ;
        RECT  1.395 6.300 13.320 6.660 ;
        RECT  8.550 6.255 9.000 6.705 ;
        RECT  4.320 6.255 4.770 6.705 ;
        RECT  1.395 6.255 1.845 6.705 ;
        LAYER metal1 ;
        RECT  12.870 6.255 13.320 6.705 ;
        RECT  8.550 6.255 9.000 6.705 ;
        RECT  4.320 6.255 4.770 6.705 ;
        RECT  1.395 6.255 1.845 6.705 ;
        END
    END a
    PIN co
        DIRECTION OUTPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  7.470 3.870 8.325 4.230 ;
        RECT  7.470 2.160 7.830 9.270 ;
        END
    END co
    PIN s
        DIRECTION OUTPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  16.830 2.160 17.190 9.270 ;
        END
    END s
    PIN ci
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  14.715 4.725 14.985 4.995 ;
        RECT  10.125 4.725 10.395 4.995 ;
        RECT  3.915 4.725 4.185 4.995 ;
        LAYER metal2 ;
        RECT  14.625 4.635 15.075 5.085 ;
        RECT  3.825 4.680 15.075 5.040 ;
        RECT  10.035 4.635 10.485 5.085 ;
        RECT  3.825 4.635 4.275 5.085 ;
        LAYER metal1 ;
        RECT  14.625 4.635 15.075 5.085 ;
        RECT  10.035 4.635 10.485 5.085 ;
        RECT  3.825 4.635 4.275 5.085 ;
        END
    END ci
    PIN b
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  13.500 5.535 13.770 5.805 ;
        RECT  9.360 5.535 9.630 5.805 ;
        RECT  5.940 5.535 6.210 5.805 ;
        RECT  2.295 5.535 2.565 5.805 ;
        LAYER metal2 ;
        RECT  13.410 5.445 13.860 5.895 ;
        RECT  2.115 5.490 13.860 5.850 ;
        RECT  9.270 5.445 9.720 5.895 ;
        RECT  5.850 5.445 6.300 5.895 ;
        RECT  2.205 5.445 2.655 5.895 ;
        LAYER metal1 ;
        RECT  13.410 5.445 13.860 5.895 ;
        RECT  9.270 5.445 9.720 5.895 ;
        RECT  5.850 5.445 6.300 5.895 ;
        RECT  2.205 5.445 2.655 5.895 ;
        END
    END b
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 17.820 11.340 ;
        RECT  15.885 8.010 16.245 11.340 ;
        RECT  9.720 8.010 10.080 11.340 ;
        RECT  8.235 8.010 8.595 11.340 ;
        RECT  6.660 8.010 7.020 11.340 ;
        RECT  2.160 8.010 2.520 11.340 ;
        RECT  0.630 8.010 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 17.820 0.990 ;
        RECT  15.840 0.000 16.200 2.790 ;
        RECT  15.030 0.000 15.390 2.790 ;
        RECT  13.500 0.000 13.860 2.790 ;
        RECT  8.190 0.000 8.550 2.790 ;
        RECT  6.705 0.000 7.065 2.790 ;
        RECT  5.985 0.000 6.345 2.790 ;
        RECT  4.365 0.000 4.725 2.790 ;
        RECT  0.630 0.000 0.990 2.655 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  1.350 8.685 1.800 9.135 ;
        RECT  1.395 8.010 1.755 9.270 ;
        RECT  3.600 2.205 4.050 2.655 ;
        RECT  3.600 8.685 4.050 9.135 ;
        RECT  3.600 8.775 4.770 9.135 ;
        RECT  3.645 8.010 4.005 9.270 ;
        RECT  4.410 8.010 4.770 9.270 ;
        RECT  5.085 2.205 5.535 2.655 ;
        RECT  2.160 2.295 3.240 2.655 ;
        RECT  2.880 2.295 3.240 4.230 ;
        RECT  2.880 3.870 5.535 4.230 ;
        RECT  5.175 3.870 5.535 7.470 ;
        RECT  2.880 7.110 6.570 7.470 ;
        RECT  6.120 7.065 6.570 7.515 ;
        RECT  2.880 7.110 3.240 9.270 ;
        RECT  5.895 7.110 6.255 9.270 ;
        RECT  8.910 8.685 9.360 9.135 ;
        RECT  8.955 8.010 9.315 9.270 ;
        RECT  10.395 8.685 10.845 9.135 ;
        RECT  10.440 8.010 10.800 9.270 ;
        RECT  12.510 7.065 12.960 7.515 ;
        RECT  11.925 8.010 12.285 9.270 ;
        RECT  11.880 8.685 12.330 9.135 ;
        RECT  12.735 8.010 13.095 9.270 ;
        RECT  11.925 8.910 13.095 9.270 ;
        RECT  12.735 2.205 13.185 2.655 ;
        RECT  11.970 2.295 13.185 2.655 ;
        RECT  14.220 2.205 14.670 2.655 ;
        RECT  10.485 2.295 11.565 2.655 ;
        RECT  11.205 3.870 16.065 4.230 ;
        RECT  15.705 3.870 16.065 7.470 ;
        RECT  15.030 7.110 16.065 7.470 ;
        RECT  11.205 2.295 11.565 9.270 ;
        RECT  15.030 7.110 15.390 9.270 ;
        LAYER via ;
        RECT  1.440 8.775 1.710 9.045 ;
        RECT  3.690 8.775 3.960 9.045 ;
        RECT  3.690 2.295 3.960 2.565 ;
        RECT  5.175 2.295 5.445 2.565 ;
        RECT  6.210 7.155 6.480 7.425 ;
        RECT  9.000 8.775 9.270 9.045 ;
        RECT  10.485 8.775 10.755 9.045 ;
        RECT  11.970 8.775 12.240 9.045 ;
        RECT  12.600 7.155 12.870 7.425 ;
        RECT  12.825 2.295 13.095 2.565 ;
        RECT  14.310 2.295 14.580 2.565 ;
        LAYER metal2 ;
        RECT  1.350 8.730 4.095 9.090 ;
        RECT  1.350 8.685 1.800 9.135 ;
        RECT  3.600 8.685 4.050 9.135 ;
        RECT  3.600 2.250 5.535 2.610 ;
        RECT  3.600 2.205 4.050 2.655 ;
        RECT  5.085 2.205 5.535 2.655 ;
        RECT  8.910 8.730 12.330 9.090 ;
        RECT  8.910 8.685 9.360 9.135 ;
        RECT  10.395 8.685 10.845 9.135 ;
        RECT  11.880 8.685 12.330 9.135 ;
        RECT  6.120 7.110 12.960 7.470 ;
        RECT  6.120 7.065 6.570 7.515 ;
        RECT  12.510 7.065 12.960 7.515 ;
        RECT  12.735 2.250 14.670 2.610 ;
        RECT  12.735 2.205 13.185 2.655 ;
        RECT  14.220 2.205 14.670 2.655 ;
    END
END fulladder

MACRO filler
    CLASS CORE ;
    FOREIGN filler 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.810 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 0.810 0.990 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 0.810 11.340 ;
        END
    END vdd!
END filler

MACRO dtrsp_2
    CLASS CORE ;
    FOREIGN dtrsp_2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 32.400 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN s
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  27.405 3.915 27.675 4.185 ;
        RECT  16.875 3.915 17.145 4.185 ;
        RECT  9.585 3.960 9.855 4.230 ;
        LAYER metal2 ;
        RECT  27.315 3.825 27.765 4.275 ;
        RECT  24.165 4.680 27.720 5.040 ;
        RECT  27.360 3.825 27.720 5.040 ;
        RECT  24.165 3.870 24.525 5.040 ;
        RECT  9.495 3.870 24.525 4.230 ;
        RECT  16.785 3.825 17.235 4.275 ;
        RECT  9.495 3.870 9.945 4.320 ;
        LAYER metal1 ;
        RECT  27.315 3.825 27.765 4.275 ;
        RECT  16.785 3.825 17.235 4.275 ;
        RECT  9.495 3.870 9.945 4.320 ;
        END
    END s
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER metal1 ;
        RECT  11.970 4.680 12.330 5.040 ;
        END
    END ck
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  4.680 5.490 5.040 5.850 ;
        END
    END ip
    PIN sm
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  5.535 6.345 5.805 6.615 ;
        RECT  1.485 6.345 1.755 6.615 ;
        LAYER metal2 ;
        RECT  5.445 6.255 5.895 6.705 ;
        RECT  1.395 6.300 5.895 6.660 ;
        RECT  1.395 6.255 1.845 6.705 ;
        LAYER metal1 ;
        RECT  5.445 6.255 5.895 6.705 ;
        RECT  1.395 6.255 1.845 6.705 ;
        END
    END sm
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  30.600 4.680 30.960 6.885 ;
        RECT  30.240 6.480 30.600 9.270 ;
        RECT  28.980 4.680 30.960 5.040 ;
        RECT  29.745 2.295 30.510 2.655 ;
        RECT  29.745 2.295 30.105 5.040 ;
        END
    END q
    PIN sip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  3.060 4.680 3.420 5.040 ;
        END
    END sip
    PIN rb
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  25.785 7.155 26.055 7.425 ;
        RECT  17.685 7.155 17.955 7.425 ;
        RECT  10.395 7.155 10.665 7.425 ;
        LAYER metal2 ;
        RECT  25.695 7.065 26.145 7.515 ;
        RECT  10.305 7.110 26.145 7.470 ;
        RECT  17.595 7.065 18.045 7.515 ;
        RECT  10.305 7.065 10.755 7.515 ;
        LAYER metal1 ;
        RECT  25.695 7.065 26.145 7.515 ;
        RECT  17.595 7.065 18.045 7.515 ;
        RECT  10.305 7.065 10.755 7.515 ;
        END
    END rb
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 32.400 11.340 ;
        RECT  31.185 8.010 31.545 11.340 ;
        RECT  29.070 8.010 29.430 11.340 ;
        RECT  25.425 8.010 25.785 11.340 ;
        RECT  22.095 8.010 22.455 11.340 ;
        RECT  19.935 8.010 20.295 11.340 ;
        RECT  17.145 8.010 17.505 11.340 ;
        RECT  11.700 8.010 12.060 11.340 ;
        RECT  10.710 8.010 11.070 11.340 ;
        RECT  8.280 8.010 8.640 11.340 ;
        RECT  6.075 8.010 6.435 11.340 ;
        RECT  1.935 8.010 2.295 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 32.400 0.990 ;
        RECT  31.140 0.000 31.500 2.655 ;
        RECT  29.070 0.000 29.430 2.655 ;
        RECT  27.360 0.000 27.720 2.655 ;
        RECT  22.095 0.000 22.455 2.655 ;
        RECT  20.115 0.000 20.475 2.655 ;
        RECT  17.505 0.000 17.865 2.655 ;
        RECT  11.745 0.000 12.105 2.655 ;
        RECT  9.090 0.000 9.450 2.655 ;
        RECT  5.850 0.000 6.210 2.655 ;
        RECT  1.890 0.000 2.250 2.655 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  0.630 3.870 2.655 4.230 ;
        RECT  2.205 3.825 2.655 4.275 ;
        RECT  0.630 2.295 0.990 9.270 ;
        RECT  5.445 3.825 5.895 4.275 ;
        RECT  3.960 4.680 7.020 5.040 ;
        RECT  3.960 2.295 4.320 9.270 ;
        RECT  7.110 2.160 7.470 4.230 ;
        RECT  7.110 3.870 8.280 4.230 ;
        RECT  7.920 4.680 9.090 5.040 ;
        RECT  7.920 3.870 8.280 6.885 ;
        RECT  7.110 6.525 8.280 6.885 ;
        RECT  7.110 6.525 7.470 9.270 ;
        RECT  8.280 2.295 8.640 3.420 ;
        RECT  9.855 2.295 10.215 3.420 ;
        RECT  8.280 3.060 10.215 3.420 ;
        RECT  9.810 8.685 10.260 9.135 ;
        RECT  9.855 8.010 10.215 9.270 ;
        RECT  10.800 2.250 11.250 2.700 ;
        RECT  11.925 6.255 12.375 6.705 ;
        RECT  11.925 3.015 12.375 3.465 ;
        RECT  12.735 4.635 13.185 5.085 ;
        RECT  12.780 2.295 13.140 9.270 ;
        RECT  13.635 8.685 14.085 9.135 ;
        RECT  13.680 8.010 14.040 9.270 ;
        RECT  13.680 2.250 14.130 2.700 ;
        RECT  15.435 8.685 15.885 9.135 ;
        RECT  15.480 8.010 15.840 9.270 ;
        RECT  15.615 2.250 16.065 2.700 ;
        RECT  15.975 3.060 16.425 3.510 ;
        RECT  16.785 5.445 17.235 5.895 ;
        RECT  18.135 8.685 18.585 9.135 ;
        RECT  18.180 8.010 18.540 9.270 ;
        RECT  16.740 2.295 17.100 3.420 ;
        RECT  18.315 2.295 18.675 3.420 ;
        RECT  16.740 3.060 18.675 3.420 ;
        RECT  19.215 2.250 19.665 2.700 ;
        RECT  17.640 5.490 20.835 5.850 ;
        RECT  17.640 5.490 18.000 6.660 ;
        RECT  14.535 6.300 18.000 6.660 ;
        RECT  14.535 2.295 14.895 9.270 ;
        RECT  21.105 5.490 22.860 5.850 ;
        RECT  21.105 5.445 21.555 5.895 ;
        RECT  21.150 2.295 21.510 9.270 ;
        RECT  23.265 3.015 23.715 3.465 ;
        RECT  23.310 3.015 23.670 5.085 ;
        RECT  23.265 4.635 23.715 5.085 ;
        RECT  22.950 2.295 24.210 2.655 ;
        RECT  24.615 8.685 25.065 9.135 ;
        RECT  24.660 8.010 25.020 9.270 ;
        RECT  24.885 6.255 25.335 6.705 ;
        RECT  25.560 3.420 26.010 3.870 ;
        RECT  27.315 8.685 27.765 9.135 ;
        RECT  27.360 8.010 27.720 9.270 ;
        RECT  26.595 2.295 26.955 3.420 ;
        RECT  28.170 2.295 28.530 3.420 ;
        RECT  26.595 3.060 28.530 3.420 ;
        RECT  24.930 2.115 25.290 5.850 ;
        RECT  23.805 5.490 30.105 5.850 ;
        RECT  29.655 5.445 30.105 5.895 ;
        RECT  23.805 5.490 24.165 9.270 ;
        RECT  30.555 3.825 31.005 4.275 ;
        LAYER via ;
        RECT  2.295 3.915 2.565 4.185 ;
        RECT  5.535 3.915 5.805 4.185 ;
        RECT  9.900 8.775 10.170 9.045 ;
        RECT  10.890 2.340 11.160 2.610 ;
        RECT  12.015 6.345 12.285 6.615 ;
        RECT  12.015 3.105 12.285 3.375 ;
        RECT  12.825 4.725 13.095 4.995 ;
        RECT  13.725 8.775 13.995 9.045 ;
        RECT  13.770 2.340 14.040 2.610 ;
        RECT  15.525 8.775 15.795 9.045 ;
        RECT  15.705 2.340 15.975 2.610 ;
        RECT  16.065 3.150 16.335 3.420 ;
        RECT  16.875 5.535 17.145 5.805 ;
        RECT  18.225 8.775 18.495 9.045 ;
        RECT  19.305 2.340 19.575 2.610 ;
        RECT  21.195 5.535 21.465 5.805 ;
        RECT  23.355 4.725 23.625 4.995 ;
        RECT  23.355 3.105 23.625 3.375 ;
        RECT  24.705 8.775 24.975 9.045 ;
        RECT  24.975 6.345 25.245 6.615 ;
        RECT  25.650 3.510 25.920 3.780 ;
        RECT  27.405 8.775 27.675 9.045 ;
        RECT  29.745 5.535 30.015 5.805 ;
        RECT  30.645 3.915 30.915 4.185 ;
        LAYER metal2 ;
        RECT  2.205 3.870 5.895 4.230 ;
        RECT  2.205 3.825 2.655 4.275 ;
        RECT  5.445 3.825 5.895 4.275 ;
        RECT  9.810 8.730 14.085 9.090 ;
        RECT  9.810 8.685 10.260 9.135 ;
        RECT  13.635 8.685 14.085 9.135 ;
        RECT  10.800 2.295 14.130 2.655 ;
        RECT  10.800 2.250 11.250 2.700 ;
        RECT  13.680 2.250 14.130 2.700 ;
        RECT  11.925 3.015 12.375 3.465 ;
        RECT  11.925 3.105 16.425 3.465 ;
        RECT  15.975 3.060 16.425 3.510 ;
        RECT  15.435 8.730 18.585 9.090 ;
        RECT  15.435 8.685 15.885 9.135 ;
        RECT  18.135 8.685 18.585 9.135 ;
        RECT  15.615 2.295 19.665 2.655 ;
        RECT  15.615 2.250 16.065 2.700 ;
        RECT  19.215 2.250 19.665 2.700 ;
        RECT  16.785 5.490 21.555 5.850 ;
        RECT  16.785 5.445 17.235 5.895 ;
        RECT  21.105 5.445 21.555 5.895 ;
        RECT  12.735 4.680 23.715 5.040 ;
        RECT  12.735 4.635 13.185 5.085 ;
        RECT  23.265 4.635 23.715 5.085 ;
        RECT  11.925 6.300 25.335 6.660 ;
        RECT  11.925 6.255 12.375 6.705 ;
        RECT  24.885 6.255 25.335 6.705 ;
        RECT  23.265 3.060 25.290 3.420 ;
        RECT  23.265 3.015 23.715 3.465 ;
        RECT  24.930 3.420 26.010 3.780 ;
        RECT  25.560 3.420 26.010 3.870 ;
        RECT  24.615 8.730 27.765 9.090 ;
        RECT  24.615 8.685 25.065 9.135 ;
        RECT  27.315 8.685 27.765 9.135 ;
        RECT  29.700 3.870 31.005 4.230 ;
        RECT  30.555 3.825 31.005 4.275 ;
        RECT  29.700 3.870 30.060 5.895 ;
        RECT  29.655 5.445 30.105 5.895 ;
    END
END dtrsp_2

MACRO drsp_4
    CLASS CORE ;
    FOREIGN drsp_4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.060 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  18.540 4.680 19.935 5.040 ;
        RECT  19.575 2.160 19.935 5.040 ;
        RECT  19.260 4.680 19.620 6.660 ;
        RECT  19.080 6.210 19.440 9.270 ;
        END
    END q
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER metal1 ;
        RECT  3.870 4.680 4.230 5.040 ;
        END
    END ck
    PIN s
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  16.875 4.725 17.145 4.995 ;
        RECT  7.245 3.915 7.515 4.185 ;
        RECT  1.485 3.915 1.755 4.185 ;
        LAYER metal2 ;
        RECT  16.785 4.635 17.235 5.085 ;
        RECT  14.490 4.680 17.235 5.040 ;
        RECT  14.490 3.870 14.850 5.040 ;
        RECT  1.395 3.870 14.850 4.230 ;
        RECT  7.155 3.825 7.605 4.275 ;
        RECT  1.395 3.825 1.845 4.275 ;
        LAYER metal1 ;
        RECT  16.785 4.635 17.235 5.085 ;
        RECT  7.155 3.825 7.605 4.275 ;
        RECT  1.395 3.825 1.845 4.275 ;
        END
    END s
    PIN rb
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  15.300 7.155 15.570 7.425 ;
        RECT  8.865 7.155 9.135 7.425 ;
        RECT  2.295 7.155 2.565 7.425 ;
        LAYER metal2 ;
        RECT  15.210 7.065 15.660 7.515 ;
        RECT  2.205 7.110 15.660 7.470 ;
        RECT  8.775 7.065 9.225 7.515 ;
        RECT  2.205 7.065 2.655 7.515 ;
        LAYER metal1 ;
        RECT  15.210 7.065 15.660 7.515 ;
        RECT  8.775 7.065 9.225 7.515 ;
        RECT  2.205 7.065 2.655 7.515 ;
        END
    END rb
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 21.060 11.340 ;
        RECT  19.890 6.750 20.250 11.340 ;
        RECT  18.315 6.750 18.675 11.340 ;
        RECT  15.660 8.010 16.020 11.340 ;
        RECT  12.690 8.010 13.050 11.340 ;
        RECT  11.115 8.010 11.475 11.340 ;
        RECT  8.190 8.010 8.550 11.340 ;
        RECT  3.465 8.010 3.825 11.340 ;
        RECT  2.655 8.010 3.015 11.340 ;
        RECT  0.630 8.010 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 21.060 0.990 ;
        RECT  20.340 0.000 20.700 3.420 ;
        RECT  18.810 0.000 19.170 3.420 ;
        RECT  17.280 0.000 17.640 3.420 ;
        RECT  12.960 0.000 13.320 2.790 ;
        RECT  11.340 0.000 11.700 2.790 ;
        RECT  8.955 0.000 9.315 2.790 ;
        RECT  3.780 0.000 4.140 2.655 ;
        RECT  1.350 0.000 1.710 2.790 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  1.890 8.685 2.340 9.135 ;
        RECT  1.935 8.010 2.295 9.270 ;
        RECT  0.630 2.160 0.990 3.420 ;
        RECT  2.115 2.160 2.475 3.420 ;
        RECT  0.630 3.060 2.475 3.420 ;
        RECT  2.790 2.205 3.240 2.655 ;
        RECT  3.465 3.015 3.915 3.465 ;
        RECT  3.735 6.255 4.185 6.705 ;
        RECT  4.500 4.635 4.950 5.085 ;
        RECT  4.545 2.160 4.905 7.560 ;
        RECT  4.230 7.200 4.590 9.270 ;
        RECT  5.220 8.685 5.670 9.135 ;
        RECT  5.265 8.010 5.625 9.270 ;
        RECT  5.355 2.205 5.805 2.655 ;
        RECT  6.750 8.685 7.200 9.135 ;
        RECT  6.795 8.010 7.155 9.270 ;
        RECT  6.885 2.205 7.335 2.655 ;
        RECT  7.065 3.015 7.515 3.465 ;
        RECT  8.910 8.685 9.360 9.135 ;
        RECT  8.955 8.010 9.315 9.270 ;
        RECT  9.270 5.445 9.720 5.895 ;
        RECT  8.235 2.160 8.595 3.420 ;
        RECT  9.720 2.160 10.080 3.420 ;
        RECT  8.235 3.060 10.080 3.420 ;
        RECT  10.440 2.205 10.890 2.655 ;
        RECT  6.165 2.160 6.525 5.850 ;
        RECT  10.350 5.490 11.565 5.850 ;
        RECT  10.350 5.490 10.710 6.660 ;
        RECT  6.030 6.300 10.710 6.660 ;
        RECT  6.030 5.490 6.390 9.270 ;
        RECT  12.105 2.160 12.465 5.850 ;
        RECT  11.925 5.445 12.465 5.850 ;
        RECT  11.880 5.490 13.140 5.850 ;
        RECT  11.880 5.490 12.375 5.895 ;
        RECT  11.880 5.490 12.240 9.270 ;
        RECT  13.905 3.015 14.355 3.465 ;
        RECT  13.680 3.420 14.310 3.780 ;
        RECT  13.680 3.420 14.040 5.085 ;
        RECT  13.635 4.635 14.085 5.085 ;
        RECT  13.725 2.295 14.805 2.655 ;
        RECT  14.445 6.255 14.895 6.705 ;
        RECT  14.850 8.685 15.300 9.135 ;
        RECT  14.895 8.010 15.255 9.270 ;
        RECT  15.435 3.825 15.885 4.275 ;
        RECT  16.920 8.685 17.370 9.135 ;
        RECT  16.965 6.750 17.325 9.270 ;
        RECT  16.560 2.160 16.920 4.230 ;
        RECT  18.045 2.160 18.405 4.230 ;
        RECT  16.560 3.870 18.405 4.230 ;
        RECT  15.210 2.160 15.570 3.420 ;
        RECT  14.715 3.060 15.570 3.420 ;
        RECT  14.715 3.060 15.075 5.850 ;
        RECT  13.590 5.490 18.900 5.850 ;
        RECT  13.590 5.490 13.950 7.470 ;
        RECT  13.590 7.110 14.445 7.470 ;
        RECT  14.085 7.110 14.445 9.270 ;
        LAYER via ;
        RECT  1.980 8.775 2.250 9.045 ;
        RECT  2.880 2.295 3.150 2.565 ;
        RECT  3.555 3.105 3.825 3.375 ;
        RECT  3.825 6.345 4.095 6.615 ;
        RECT  4.590 4.725 4.860 4.995 ;
        RECT  5.310 8.775 5.580 9.045 ;
        RECT  5.445 2.295 5.715 2.565 ;
        RECT  6.840 8.775 7.110 9.045 ;
        RECT  6.975 2.295 7.245 2.565 ;
        RECT  7.155 3.105 7.425 3.375 ;
        RECT  9.000 8.775 9.270 9.045 ;
        RECT  9.360 5.535 9.630 5.805 ;
        RECT  10.530 2.295 10.800 2.565 ;
        RECT  12.015 5.535 12.285 5.805 ;
        RECT  13.725 4.725 13.995 4.995 ;
        RECT  13.995 3.105 14.265 3.375 ;
        RECT  14.535 6.345 14.805 6.615 ;
        RECT  14.940 8.775 15.210 9.045 ;
        RECT  15.525 3.915 15.795 4.185 ;
        RECT  17.010 8.775 17.280 9.045 ;
        LAYER metal2 ;
        RECT  1.890 8.730 5.670 9.090 ;
        RECT  1.890 8.685 2.340 9.135 ;
        RECT  5.220 8.685 5.670 9.135 ;
        RECT  2.790 2.250 5.805 2.610 ;
        RECT  2.790 2.205 3.240 2.655 ;
        RECT  5.355 2.205 5.805 2.655 ;
        RECT  3.465 3.060 7.515 3.420 ;
        RECT  3.465 3.015 3.915 3.465 ;
        RECT  7.065 3.015 7.515 3.465 ;
        RECT  6.750 8.730 9.360 9.090 ;
        RECT  6.750 8.685 7.200 9.135 ;
        RECT  8.910 8.685 9.360 9.135 ;
        RECT  6.885 2.250 10.890 2.610 ;
        RECT  6.885 2.205 7.335 2.655 ;
        RECT  10.440 2.205 10.890 2.655 ;
        RECT  9.270 5.490 12.375 5.850 ;
        RECT  9.270 5.445 9.720 5.895 ;
        RECT  11.925 5.445 12.375 5.895 ;
        RECT  4.500 4.680 14.085 5.040 ;
        RECT  4.500 4.635 4.950 5.085 ;
        RECT  13.635 4.635 14.085 5.085 ;
        RECT  3.735 6.300 14.895 6.660 ;
        RECT  3.735 6.255 4.185 6.705 ;
        RECT  14.445 6.255 14.895 6.705 ;
        RECT  13.905 3.060 15.570 3.420 ;
        RECT  13.905 3.015 14.355 3.465 ;
        RECT  15.210 3.060 15.570 4.230 ;
        RECT  15.435 3.825 15.885 4.275 ;
        RECT  14.850 8.730 17.370 9.090 ;
        RECT  14.850 8.685 15.300 9.135 ;
        RECT  16.920 8.685 17.370 9.135 ;
    END
END drsp_4

MACRO drsp_2
    CLASS CORE ;
    FOREIGN drsp_2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.060 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  19.080 6.750 20.430 7.110 ;
        RECT  20.070 4.680 20.430 7.110 ;
        RECT  18.540 4.680 20.430 5.040 ;
        RECT  19.575 2.160 19.935 5.040 ;
        RECT  19.080 6.750 19.440 9.270 ;
        END
    END q
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER metal1 ;
        RECT  3.870 4.680 4.230 5.040 ;
        END
    END ck
    PIN s
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  16.875 4.725 17.145 4.995 ;
        RECT  7.245 3.915 7.515 4.185 ;
        RECT  1.485 3.915 1.755 4.185 ;
        LAYER metal2 ;
        RECT  16.785 4.635 17.235 5.085 ;
        RECT  14.490 4.680 17.235 5.040 ;
        RECT  14.490 3.870 14.850 5.040 ;
        RECT  1.395 3.870 14.850 4.230 ;
        RECT  7.155 3.825 7.605 4.275 ;
        RECT  1.395 3.825 1.845 4.275 ;
        LAYER metal1 ;
        RECT  16.785 4.635 17.235 5.085 ;
        RECT  7.155 3.825 7.605 4.275 ;
        RECT  1.395 3.825 1.845 4.275 ;
        END
    END s
    PIN rb
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  15.300 7.155 15.570 7.425 ;
        RECT  8.865 7.155 9.135 7.425 ;
        RECT  2.295 7.155 2.565 7.425 ;
        LAYER metal2 ;
        RECT  15.210 7.065 15.660 7.515 ;
        RECT  2.205 7.110 15.660 7.470 ;
        RECT  8.775 7.065 9.225 7.515 ;
        RECT  2.205 7.065 2.655 7.515 ;
        LAYER metal1 ;
        RECT  15.210 7.065 15.660 7.515 ;
        RECT  8.775 7.065 9.225 7.515 ;
        RECT  2.205 7.065 2.655 7.515 ;
        END
    END rb
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 21.060 11.340 ;
        RECT  18.315 6.750 18.675 11.340 ;
        RECT  15.660 8.010 16.020 11.340 ;
        RECT  12.690 8.010 13.050 11.340 ;
        RECT  11.115 8.010 11.475 11.340 ;
        RECT  8.190 8.010 8.550 11.340 ;
        RECT  3.465 8.010 3.825 11.340 ;
        RECT  2.655 8.010 3.015 11.340 ;
        RECT  0.630 8.010 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 21.060 0.990 ;
        RECT  18.810 0.000 19.170 3.420 ;
        RECT  17.280 0.000 17.640 3.420 ;
        RECT  12.960 0.000 13.320 2.790 ;
        RECT  11.340 0.000 11.700 2.790 ;
        RECT  8.955 0.000 9.315 2.790 ;
        RECT  3.780 0.000 4.140 2.655 ;
        RECT  1.350 0.000 1.710 2.790 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  1.890 8.685 2.340 9.135 ;
        RECT  1.935 8.010 2.295 9.270 ;
        RECT  0.630 2.160 0.990 3.420 ;
        RECT  2.115 2.160 2.475 3.420 ;
        RECT  0.630 3.060 2.475 3.420 ;
        RECT  2.790 2.205 3.240 2.655 ;
        RECT  3.465 3.015 3.915 3.465 ;
        RECT  3.735 6.255 4.185 6.705 ;
        RECT  4.500 4.635 4.950 5.085 ;
        RECT  4.545 2.160 4.905 7.560 ;
        RECT  4.230 7.200 4.590 9.270 ;
        RECT  5.220 8.685 5.670 9.135 ;
        RECT  5.265 8.010 5.625 9.270 ;
        RECT  5.355 2.205 5.805 2.655 ;
        RECT  6.750 8.685 7.200 9.135 ;
        RECT  6.795 8.010 7.155 9.270 ;
        RECT  6.885 2.205 7.335 2.655 ;
        RECT  7.065 3.015 7.515 3.465 ;
        RECT  8.910 8.685 9.360 9.135 ;
        RECT  8.955 8.010 9.315 9.270 ;
        RECT  9.270 5.445 9.720 5.895 ;
        RECT  8.235 2.160 8.595 3.420 ;
        RECT  9.720 2.160 10.080 3.420 ;
        RECT  8.235 3.060 10.080 3.420 ;
        RECT  10.440 2.205 10.890 2.655 ;
        RECT  6.165 2.160 6.525 5.850 ;
        RECT  10.350 5.490 11.565 5.850 ;
        RECT  10.350 5.490 10.710 6.660 ;
        RECT  6.030 6.300 10.710 6.660 ;
        RECT  6.030 5.490 6.390 9.270 ;
        RECT  12.105 2.160 12.465 5.850 ;
        RECT  11.925 5.445 12.465 5.850 ;
        RECT  11.880 5.490 13.140 5.850 ;
        RECT  11.880 5.490 12.375 5.895 ;
        RECT  11.880 5.490 12.240 9.270 ;
        RECT  13.905 3.015 14.355 3.465 ;
        RECT  13.680 3.420 14.310 3.780 ;
        RECT  13.680 3.420 14.040 5.085 ;
        RECT  13.635 4.635 14.085 5.085 ;
        RECT  13.725 2.295 14.805 2.655 ;
        RECT  14.445 6.255 14.895 6.705 ;
        RECT  14.850 8.685 15.300 9.135 ;
        RECT  14.895 8.010 15.255 9.270 ;
        RECT  15.435 3.825 15.885 4.275 ;
        RECT  16.920 8.685 17.370 9.135 ;
        RECT  16.965 6.750 17.325 9.270 ;
        RECT  16.560 2.160 16.920 4.230 ;
        RECT  18.045 2.160 18.405 4.230 ;
        RECT  16.560 3.870 18.405 4.230 ;
        RECT  15.210 2.160 15.570 3.420 ;
        RECT  14.715 3.060 15.570 3.420 ;
        RECT  14.715 3.060 15.075 5.850 ;
        RECT  13.590 5.490 18.990 5.850 ;
        RECT  13.590 5.490 13.950 7.470 ;
        RECT  13.590 7.110 14.445 7.470 ;
        RECT  14.085 7.110 14.445 9.270 ;
        LAYER via ;
        RECT  1.980 8.775 2.250 9.045 ;
        RECT  2.880 2.295 3.150 2.565 ;
        RECT  3.555 3.105 3.825 3.375 ;
        RECT  3.825 6.345 4.095 6.615 ;
        RECT  4.590 4.725 4.860 4.995 ;
        RECT  5.310 8.775 5.580 9.045 ;
        RECT  5.445 2.295 5.715 2.565 ;
        RECT  6.840 8.775 7.110 9.045 ;
        RECT  6.975 2.295 7.245 2.565 ;
        RECT  7.155 3.105 7.425 3.375 ;
        RECT  9.000 8.775 9.270 9.045 ;
        RECT  9.360 5.535 9.630 5.805 ;
        RECT  10.530 2.295 10.800 2.565 ;
        RECT  12.015 5.535 12.285 5.805 ;
        RECT  13.725 4.725 13.995 4.995 ;
        RECT  13.995 3.105 14.265 3.375 ;
        RECT  14.535 6.345 14.805 6.615 ;
        RECT  14.940 8.775 15.210 9.045 ;
        RECT  15.525 3.915 15.795 4.185 ;
        RECT  17.010 8.775 17.280 9.045 ;
        LAYER metal2 ;
        RECT  1.890 8.730 5.670 9.090 ;
        RECT  1.890 8.685 2.340 9.135 ;
        RECT  5.220 8.685 5.670 9.135 ;
        RECT  2.790 2.250 5.805 2.610 ;
        RECT  2.790 2.205 3.240 2.655 ;
        RECT  5.355 2.205 5.805 2.655 ;
        RECT  3.465 3.060 7.515 3.420 ;
        RECT  3.465 3.015 3.915 3.465 ;
        RECT  7.065 3.015 7.515 3.465 ;
        RECT  6.750 8.730 9.360 9.090 ;
        RECT  6.750 8.685 7.200 9.135 ;
        RECT  8.910 8.685 9.360 9.135 ;
        RECT  6.885 2.250 10.890 2.610 ;
        RECT  6.885 2.205 7.335 2.655 ;
        RECT  10.440 2.205 10.890 2.655 ;
        RECT  9.270 5.490 12.375 5.850 ;
        RECT  9.270 5.445 9.720 5.895 ;
        RECT  11.925 5.445 12.375 5.895 ;
        RECT  4.500 4.680 14.085 5.040 ;
        RECT  4.500 4.635 4.950 5.085 ;
        RECT  13.635 4.635 14.085 5.085 ;
        RECT  3.735 6.300 14.895 6.660 ;
        RECT  3.735 6.255 4.185 6.705 ;
        RECT  14.445 6.255 14.895 6.705 ;
        RECT  13.905 3.060 15.570 3.420 ;
        RECT  13.905 3.015 14.355 3.465 ;
        RECT  15.210 3.060 15.570 4.230 ;
        RECT  15.435 3.825 15.885 4.275 ;
        RECT  14.850 8.730 17.370 9.090 ;
        RECT  14.850 8.685 15.300 9.135 ;
        RECT  16.920 8.685 17.370 9.135 ;
    END
END drsp_2

MACRO drsp_1
    CLASS CORE ;
    FOREIGN drsp_1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.060 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip
    PIN rb
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  15.300 7.155 15.570 7.425 ;
        RECT  8.865 7.155 9.135 7.425 ;
        RECT  2.295 7.155 2.565 7.425 ;
        LAYER metal2 ;
        RECT  15.210 7.065 15.660 7.515 ;
        RECT  2.205 7.110 15.660 7.470 ;
        RECT  8.775 7.065 9.225 7.515 ;
        RECT  2.205 7.065 2.655 7.515 ;
        LAYER metal1 ;
        RECT  15.210 7.065 15.660 7.515 ;
        RECT  8.775 7.065 9.225 7.515 ;
        RECT  2.205 7.065 2.655 7.515 ;
        END
    END rb
    PIN s
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  16.875 4.725 17.145 4.995 ;
        RECT  7.245 3.915 7.515 4.185 ;
        RECT  1.485 3.915 1.755 4.185 ;
        LAYER metal2 ;
        RECT  16.785 4.635 17.235 5.085 ;
        RECT  14.490 4.680 17.235 5.040 ;
        RECT  14.490 3.870 14.850 5.040 ;
        RECT  1.395 3.870 14.850 4.230 ;
        RECT  7.155 3.825 7.605 4.275 ;
        RECT  1.395 3.825 1.845 4.275 ;
        LAYER metal1 ;
        RECT  16.785 4.635 17.235 5.085 ;
        RECT  7.155 3.825 7.605 4.275 ;
        RECT  1.395 3.825 1.845 4.275 ;
        END
    END s
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER metal1 ;
        RECT  3.870 4.680 4.230 5.040 ;
        END
    END ck
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  19.080 6.975 20.430 7.335 ;
        RECT  20.070 4.095 20.430 7.335 ;
        RECT  18.540 4.095 20.430 4.455 ;
        RECT  19.575 2.160 19.935 4.455 ;
        RECT  19.080 6.975 19.440 9.270 ;
        END
    END q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 21.060 0.990 ;
        RECT  18.810 0.000 19.170 2.790 ;
        RECT  17.280 0.000 17.640 2.790 ;
        RECT  12.960 0.000 13.320 2.790 ;
        RECT  11.340 0.000 11.700 2.790 ;
        RECT  8.955 0.000 9.315 2.790 ;
        RECT  3.780 0.000 4.140 2.655 ;
        RECT  1.350 0.000 1.710 2.790 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 21.060 11.340 ;
        RECT  18.315 8.010 18.675 11.340 ;
        RECT  15.660 8.010 16.020 11.340 ;
        RECT  12.690 8.010 13.050 11.340 ;
        RECT  11.115 8.010 11.475 11.340 ;
        RECT  8.190 8.010 8.550 11.340 ;
        RECT  3.465 8.010 3.825 11.340 ;
        RECT  2.655 8.010 3.015 11.340 ;
        RECT  0.630 8.010 0.990 11.340 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  1.890 8.685 2.340 9.135 ;
        RECT  1.935 8.010 2.295 9.270 ;
        RECT  0.630 2.160 0.990 3.420 ;
        RECT  2.115 2.160 2.475 3.420 ;
        RECT  0.630 3.060 2.475 3.420 ;
        RECT  2.790 2.205 3.240 2.655 ;
        RECT  3.465 3.015 3.915 3.465 ;
        RECT  3.735 6.255 4.185 6.705 ;
        RECT  4.500 4.635 4.950 5.085 ;
        RECT  4.545 2.160 4.905 7.560 ;
        RECT  4.230 7.200 4.590 9.270 ;
        RECT  5.220 8.685 5.670 9.135 ;
        RECT  5.265 8.010 5.625 9.270 ;
        RECT  5.355 2.205 5.805 2.655 ;
        RECT  6.750 8.685 7.200 9.135 ;
        RECT  6.795 8.010 7.155 9.270 ;
        RECT  6.885 2.205 7.335 2.655 ;
        RECT  7.065 3.015 7.515 3.465 ;
        RECT  8.910 8.685 9.360 9.135 ;
        RECT  8.955 8.010 9.315 9.270 ;
        RECT  9.270 5.445 9.720 5.895 ;
        RECT  8.235 2.160 8.595 3.420 ;
        RECT  9.720 2.160 10.080 3.420 ;
        RECT  8.235 3.060 10.080 3.420 ;
        RECT  10.440 2.205 10.890 2.655 ;
        RECT  6.165 2.160 6.525 5.850 ;
        RECT  10.350 5.490 11.565 5.850 ;
        RECT  10.350 5.490 10.710 6.660 ;
        RECT  6.030 6.300 10.710 6.660 ;
        RECT  6.030 5.490 6.390 9.270 ;
        RECT  12.105 2.160 12.465 5.850 ;
        RECT  11.925 5.445 12.465 5.850 ;
        RECT  11.880 5.490 13.140 5.850 ;
        RECT  11.880 5.490 12.375 5.895 ;
        RECT  11.880 5.490 12.240 9.270 ;
        RECT  13.905 3.015 14.355 3.465 ;
        RECT  13.680 3.420 14.310 3.780 ;
        RECT  13.680 3.420 14.040 5.085 ;
        RECT  13.635 4.635 14.085 5.085 ;
        RECT  13.725 2.295 14.805 2.655 ;
        RECT  14.445 6.255 14.895 6.705 ;
        RECT  14.850 8.685 15.300 9.135 ;
        RECT  14.895 8.010 15.255 9.270 ;
        RECT  15.435 3.825 15.885 4.275 ;
        RECT  16.920 8.685 17.370 9.135 ;
        RECT  16.965 8.010 17.325 9.270 ;
        RECT  16.560 2.160 16.920 3.420 ;
        RECT  18.045 2.160 18.405 3.420 ;
        RECT  16.560 3.060 18.405 3.420 ;
        RECT  15.210 2.160 15.570 3.420 ;
        RECT  14.715 3.060 15.570 3.420 ;
        RECT  14.715 3.060 15.075 5.850 ;
        RECT  13.590 5.490 18.990 5.850 ;
        RECT  13.590 5.490 13.950 7.470 ;
        RECT  13.590 7.110 14.445 7.470 ;
        RECT  14.085 7.110 14.445 9.270 ;
        LAYER via ;
        RECT  1.980 8.775 2.250 9.045 ;
        RECT  2.880 2.295 3.150 2.565 ;
        RECT  3.555 3.105 3.825 3.375 ;
        RECT  3.825 6.345 4.095 6.615 ;
        RECT  4.590 4.725 4.860 4.995 ;
        RECT  5.310 8.775 5.580 9.045 ;
        RECT  5.445 2.295 5.715 2.565 ;
        RECT  6.840 8.775 7.110 9.045 ;
        RECT  6.975 2.295 7.245 2.565 ;
        RECT  7.155 3.105 7.425 3.375 ;
        RECT  9.000 8.775 9.270 9.045 ;
        RECT  9.360 5.535 9.630 5.805 ;
        RECT  10.530 2.295 10.800 2.565 ;
        RECT  12.015 5.535 12.285 5.805 ;
        RECT  13.725 4.725 13.995 4.995 ;
        RECT  13.995 3.105 14.265 3.375 ;
        RECT  14.535 6.345 14.805 6.615 ;
        RECT  14.940 8.775 15.210 9.045 ;
        RECT  15.525 3.915 15.795 4.185 ;
        RECT  17.010 8.775 17.280 9.045 ;
        LAYER metal2 ;
        RECT  1.890 8.730 5.670 9.090 ;
        RECT  1.890 8.685 2.340 9.135 ;
        RECT  5.220 8.685 5.670 9.135 ;
        RECT  2.790 2.250 5.805 2.610 ;
        RECT  2.790 2.205 3.240 2.655 ;
        RECT  5.355 2.205 5.805 2.655 ;
        RECT  3.465 3.060 7.515 3.420 ;
        RECT  3.465 3.015 3.915 3.465 ;
        RECT  7.065 3.015 7.515 3.465 ;
        RECT  6.750 8.730 9.360 9.090 ;
        RECT  6.750 8.685 7.200 9.135 ;
        RECT  8.910 8.685 9.360 9.135 ;
        RECT  6.885 2.250 10.890 2.610 ;
        RECT  6.885 2.205 7.335 2.655 ;
        RECT  10.440 2.205 10.890 2.655 ;
        RECT  9.270 5.490 12.375 5.850 ;
        RECT  9.270 5.445 9.720 5.895 ;
        RECT  11.925 5.445 12.375 5.895 ;
        RECT  4.500 4.680 14.085 5.040 ;
        RECT  4.500 4.635 4.950 5.085 ;
        RECT  13.635 4.635 14.085 5.085 ;
        RECT  3.735 6.300 14.895 6.660 ;
        RECT  3.735 6.255 4.185 6.705 ;
        RECT  14.445 6.255 14.895 6.705 ;
        RECT  13.905 3.060 15.570 3.420 ;
        RECT  13.905 3.015 14.355 3.465 ;
        RECT  15.210 3.060 15.570 4.230 ;
        RECT  15.435 3.825 15.885 4.275 ;
        RECT  14.850 8.730 17.370 9.090 ;
        RECT  14.850 8.685 15.300 9.135 ;
        RECT  16.920 8.685 17.370 9.135 ;
    END
END drsp_1

MACRO drp_4
    CLASS CORE ;
    FOREIGN drp_4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.440 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip
    PIN rb
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  14.175 7.155 14.445 7.425 ;
        RECT  7.740 7.155 8.010 7.425 ;
        RECT  1.485 7.155 1.755 7.425 ;
        LAYER metal2 ;
        RECT  14.085 7.065 14.535 7.515 ;
        RECT  1.395 7.110 14.535 7.470 ;
        RECT  7.650 7.065 8.100 7.515 ;
        RECT  1.395 7.065 1.845 7.515 ;
        LAYER metal1 ;
        RECT  14.085 7.065 14.535 7.515 ;
        RECT  7.650 7.065 8.100 7.515 ;
        RECT  1.395 7.065 1.845 7.515 ;
        END
    END rb
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER metal1 ;
        RECT  3.060 4.680 3.420 5.040 ;
        END
    END ck
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  17.370 6.120 18.810 6.480 ;
        RECT  18.450 4.095 18.810 6.480 ;
        RECT  16.830 4.095 18.810 4.455 ;
        RECT  17.865 2.160 18.225 4.455 ;
        RECT  17.370 6.120 17.730 9.270 ;
        END
    END q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 19.440 11.340 ;
        RECT  18.225 6.750 18.585 11.340 ;
        RECT  16.605 6.750 16.965 11.340 ;
        RECT  14.535 8.010 14.895 11.340 ;
        RECT  11.565 8.010 11.925 11.340 ;
        RECT  9.990 8.010 10.350 11.340 ;
        RECT  7.065 8.010 7.425 11.340 ;
        RECT  2.925 8.010 3.285 11.340 ;
        RECT  2.115 8.010 2.475 11.340 ;
        RECT  0.630 8.010 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 19.440 0.990 ;
        RECT  18.720 0.000 19.080 3.420 ;
        RECT  17.100 0.000 17.460 3.420 ;
        RECT  11.835 0.000 12.195 2.790 ;
        RECT  10.215 0.000 10.575 2.790 ;
        RECT  7.830 0.000 8.190 2.790 ;
        RECT  3.240 0.000 3.600 2.655 ;
        RECT  0.630 0.000 0.990 2.790 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  1.350 8.685 1.800 9.135 ;
        RECT  1.395 8.010 1.755 9.270 ;
        RECT  2.250 2.205 2.700 2.655 ;
        RECT  2.925 3.015 3.375 3.465 ;
        RECT  3.195 6.255 3.645 6.705 ;
        RECT  3.960 4.635 4.410 5.085 ;
        RECT  4.005 2.160 4.365 7.560 ;
        RECT  3.690 7.200 4.050 9.270 ;
        RECT  4.680 8.685 5.130 9.135 ;
        RECT  4.725 8.010 5.085 9.270 ;
        RECT  4.815 2.205 5.265 2.655 ;
        RECT  6.210 8.685 6.660 9.135 ;
        RECT  6.255 8.010 6.615 9.270 ;
        RECT  6.345 2.205 6.795 2.655 ;
        RECT  6.525 3.015 6.975 3.465 ;
        RECT  7.785 8.685 8.235 9.135 ;
        RECT  7.830 8.010 8.190 9.270 ;
        RECT  8.145 5.445 8.595 5.895 ;
        RECT  9.315 2.205 9.765 2.655 ;
        RECT  5.625 2.160 5.985 5.850 ;
        RECT  9.225 5.490 10.440 5.850 ;
        RECT  9.225 5.490 9.585 6.660 ;
        RECT  5.490 6.300 9.585 6.660 ;
        RECT  5.490 5.490 5.850 9.270 ;
        RECT  10.980 2.160 11.340 5.850 ;
        RECT  10.800 5.445 11.340 5.850 ;
        RECT  10.755 5.490 12.015 5.850 ;
        RECT  10.755 5.490 11.250 5.895 ;
        RECT  10.755 5.490 11.115 9.270 ;
        RECT  12.780 3.015 13.230 3.465 ;
        RECT  12.555 3.420 13.185 3.780 ;
        RECT  12.555 3.420 12.915 5.085 ;
        RECT  12.510 4.635 12.960 5.085 ;
        RECT  12.600 2.295 13.680 2.655 ;
        RECT  13.320 6.255 13.770 6.705 ;
        RECT  13.725 8.685 14.175 9.135 ;
        RECT  13.770 8.010 14.130 9.270 ;
        RECT  14.310 3.825 14.760 4.275 ;
        RECT  15.795 8.685 16.245 9.135 ;
        RECT  15.840 6.750 16.200 9.270 ;
        RECT  15.435 2.295 16.695 2.655 ;
        RECT  16.335 2.160 16.695 3.420 ;
        RECT  14.085 2.160 14.445 3.420 ;
        RECT  13.590 3.060 14.445 3.420 ;
        RECT  13.590 3.060 13.950 5.850 ;
        RECT  12.465 5.490 17.280 5.850 ;
        RECT  12.465 5.490 12.825 7.470 ;
        RECT  12.465 7.110 13.320 7.470 ;
        RECT  12.960 7.110 13.320 9.270 ;
        LAYER via ;
        RECT  1.440 8.775 1.710 9.045 ;
        RECT  2.340 2.295 2.610 2.565 ;
        RECT  3.015 3.105 3.285 3.375 ;
        RECT  3.285 6.345 3.555 6.615 ;
        RECT  4.050 4.725 4.320 4.995 ;
        RECT  4.770 8.775 5.040 9.045 ;
        RECT  4.905 2.295 5.175 2.565 ;
        RECT  6.300 8.775 6.570 9.045 ;
        RECT  6.435 2.295 6.705 2.565 ;
        RECT  6.615 3.105 6.885 3.375 ;
        RECT  7.875 8.775 8.145 9.045 ;
        RECT  8.235 5.535 8.505 5.805 ;
        RECT  9.405 2.295 9.675 2.565 ;
        RECT  10.890 5.535 11.160 5.805 ;
        RECT  12.600 4.725 12.870 4.995 ;
        RECT  12.870 3.105 13.140 3.375 ;
        RECT  13.410 6.345 13.680 6.615 ;
        RECT  13.815 8.775 14.085 9.045 ;
        RECT  14.400 3.915 14.670 4.185 ;
        RECT  15.885 8.775 16.155 9.045 ;
        LAYER metal2 ;
        RECT  1.350 8.730 5.130 9.090 ;
        RECT  1.350 8.685 1.800 9.135 ;
        RECT  4.680 8.685 5.130 9.135 ;
        RECT  2.250 2.250 5.265 2.610 ;
        RECT  2.250 2.205 2.700 2.655 ;
        RECT  4.815 2.205 5.265 2.655 ;
        RECT  2.925 3.060 6.975 3.420 ;
        RECT  2.925 3.015 3.375 3.465 ;
        RECT  6.525 3.015 6.975 3.465 ;
        RECT  6.210 8.730 8.235 9.090 ;
        RECT  6.210 8.685 6.660 9.135 ;
        RECT  7.785 8.685 8.235 9.135 ;
        RECT  6.345 2.250 9.765 2.610 ;
        RECT  6.345 2.205 6.795 2.655 ;
        RECT  9.315 2.205 9.765 2.655 ;
        RECT  8.145 5.490 11.250 5.850 ;
        RECT  8.145 5.445 8.595 5.895 ;
        RECT  10.800 5.445 11.250 5.895 ;
        RECT  3.960 4.680 12.960 5.040 ;
        RECT  3.960 4.635 4.410 5.085 ;
        RECT  12.510 4.635 12.960 5.085 ;
        RECT  3.195 6.300 13.770 6.660 ;
        RECT  3.195 6.255 3.645 6.705 ;
        RECT  13.320 6.255 13.770 6.705 ;
        RECT  12.780 3.060 14.445 3.420 ;
        RECT  12.780 3.015 13.230 3.465 ;
        RECT  14.085 3.060 14.445 4.230 ;
        RECT  14.310 3.825 14.760 4.275 ;
        RECT  13.725 8.730 16.245 9.090 ;
        RECT  13.725 8.685 14.175 9.135 ;
        RECT  15.795 8.685 16.245 9.135 ;
    END
END drp_4

MACRO drp_2
    CLASS CORE ;
    FOREIGN drp_2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.440 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  17.370 6.750 18.810 7.110 ;
        RECT  18.450 4.095 18.810 7.110 ;
        RECT  16.830 4.095 18.810 4.455 ;
        RECT  17.865 2.160 18.225 4.455 ;
        RECT  17.370 6.750 17.730 9.270 ;
        END
    END q
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER metal1 ;
        RECT  3.060 4.680 3.420 5.040 ;
        END
    END ck
    PIN rb
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  14.175 7.155 14.445 7.425 ;
        RECT  7.740 7.155 8.010 7.425 ;
        RECT  1.485 7.155 1.755 7.425 ;
        LAYER metal2 ;
        RECT  14.085 7.065 14.535 7.515 ;
        RECT  1.395 7.110 14.535 7.470 ;
        RECT  7.650 7.065 8.100 7.515 ;
        RECT  1.395 7.065 1.845 7.515 ;
        LAYER metal1 ;
        RECT  14.085 7.065 14.535 7.515 ;
        RECT  7.650 7.065 8.100 7.515 ;
        RECT  1.395 7.065 1.845 7.515 ;
        END
    END rb
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 19.440 11.340 ;
        RECT  16.605 6.750 16.965 11.340 ;
        RECT  14.535 8.010 14.895 11.340 ;
        RECT  11.565 8.010 11.925 11.340 ;
        RECT  9.990 8.010 10.350 11.340 ;
        RECT  7.065 8.010 7.425 11.340 ;
        RECT  2.925 8.010 3.285 11.340 ;
        RECT  2.115 8.010 2.475 11.340 ;
        RECT  0.630 8.010 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 19.440 0.990 ;
        RECT  17.100 0.000 17.460 3.420 ;
        RECT  11.835 0.000 12.195 2.790 ;
        RECT  10.215 0.000 10.575 2.790 ;
        RECT  7.830 0.000 8.190 2.790 ;
        RECT  3.240 0.000 3.600 2.655 ;
        RECT  0.630 0.000 0.990 2.790 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  1.350 8.685 1.800 9.135 ;
        RECT  1.395 8.010 1.755 9.270 ;
        RECT  2.250 2.205 2.700 2.655 ;
        RECT  2.925 3.015 3.375 3.465 ;
        RECT  3.195 6.255 3.645 6.705 ;
        RECT  3.960 4.635 4.410 5.085 ;
        RECT  4.005 2.160 4.365 7.560 ;
        RECT  3.690 7.200 4.050 9.270 ;
        RECT  4.680 8.685 5.130 9.135 ;
        RECT  4.725 8.010 5.085 9.270 ;
        RECT  4.815 2.205 5.265 2.655 ;
        RECT  6.210 8.685 6.660 9.135 ;
        RECT  6.255 8.010 6.615 9.270 ;
        RECT  6.345 2.205 6.795 2.655 ;
        RECT  6.525 3.015 6.975 3.465 ;
        RECT  7.785 8.685 8.235 9.135 ;
        RECT  7.830 8.010 8.190 9.270 ;
        RECT  8.145 5.445 8.595 5.895 ;
        RECT  9.315 2.205 9.765 2.655 ;
        RECT  5.625 2.160 5.985 5.850 ;
        RECT  9.225 5.490 10.440 5.850 ;
        RECT  9.225 5.490 9.585 6.660 ;
        RECT  5.490 6.300 9.585 6.660 ;
        RECT  5.490 5.490 5.850 9.270 ;
        RECT  10.980 2.160 11.340 5.850 ;
        RECT  10.800 5.445 11.340 5.850 ;
        RECT  10.755 5.490 12.015 5.850 ;
        RECT  10.755 5.490 11.250 5.895 ;
        RECT  10.755 5.490 11.115 9.270 ;
        RECT  12.780 3.015 13.230 3.465 ;
        RECT  12.555 3.420 13.185 3.780 ;
        RECT  12.555 3.420 12.915 5.085 ;
        RECT  12.510 4.635 12.960 5.085 ;
        RECT  12.600 2.295 13.680 2.655 ;
        RECT  13.320 6.255 13.770 6.705 ;
        RECT  13.725 8.685 14.175 9.135 ;
        RECT  13.770 8.010 14.130 9.270 ;
        RECT  14.310 3.825 14.760 4.275 ;
        RECT  15.795 8.685 16.245 9.135 ;
        RECT  15.840 6.750 16.200 9.270 ;
        RECT  15.435 2.295 16.695 2.655 ;
        RECT  16.335 2.160 16.695 3.420 ;
        RECT  14.085 2.160 14.445 3.420 ;
        RECT  13.590 3.060 14.445 3.420 ;
        RECT  13.590 3.060 13.950 5.850 ;
        RECT  12.465 5.490 17.280 5.850 ;
        RECT  12.465 5.490 12.825 7.470 ;
        RECT  12.465 7.110 13.320 7.470 ;
        RECT  12.960 7.110 13.320 9.270 ;
        LAYER via ;
        RECT  1.440 8.775 1.710 9.045 ;
        RECT  2.340 2.295 2.610 2.565 ;
        RECT  3.015 3.105 3.285 3.375 ;
        RECT  3.285 6.345 3.555 6.615 ;
        RECT  4.050 4.725 4.320 4.995 ;
        RECT  4.770 8.775 5.040 9.045 ;
        RECT  4.905 2.295 5.175 2.565 ;
        RECT  6.300 8.775 6.570 9.045 ;
        RECT  6.435 2.295 6.705 2.565 ;
        RECT  6.615 3.105 6.885 3.375 ;
        RECT  7.875 8.775 8.145 9.045 ;
        RECT  8.235 5.535 8.505 5.805 ;
        RECT  9.405 2.295 9.675 2.565 ;
        RECT  10.890 5.535 11.160 5.805 ;
        RECT  12.600 4.725 12.870 4.995 ;
        RECT  12.870 3.105 13.140 3.375 ;
        RECT  13.410 6.345 13.680 6.615 ;
        RECT  13.815 8.775 14.085 9.045 ;
        RECT  14.400 3.915 14.670 4.185 ;
        RECT  15.885 8.775 16.155 9.045 ;
        LAYER metal2 ;
        RECT  1.350 8.730 5.130 9.090 ;
        RECT  1.350 8.685 1.800 9.135 ;
        RECT  4.680 8.685 5.130 9.135 ;
        RECT  2.250 2.250 5.265 2.610 ;
        RECT  2.250 2.205 2.700 2.655 ;
        RECT  4.815 2.205 5.265 2.655 ;
        RECT  2.925 3.060 6.975 3.420 ;
        RECT  2.925 3.015 3.375 3.465 ;
        RECT  6.525 3.015 6.975 3.465 ;
        RECT  6.210 8.730 8.235 9.090 ;
        RECT  6.210 8.685 6.660 9.135 ;
        RECT  7.785 8.685 8.235 9.135 ;
        RECT  6.345 2.250 9.765 2.610 ;
        RECT  6.345 2.205 6.795 2.655 ;
        RECT  9.315 2.205 9.765 2.655 ;
        RECT  8.145 5.490 11.250 5.850 ;
        RECT  8.145 5.445 8.595 5.895 ;
        RECT  10.800 5.445 11.250 5.895 ;
        RECT  3.960 4.680 12.960 5.040 ;
        RECT  3.960 4.635 4.410 5.085 ;
        RECT  12.510 4.635 12.960 5.085 ;
        RECT  3.195 6.300 13.770 6.660 ;
        RECT  3.195 6.255 3.645 6.705 ;
        RECT  13.320 6.255 13.770 6.705 ;
        RECT  12.780 3.060 14.445 3.420 ;
        RECT  12.780 3.015 13.230 3.465 ;
        RECT  14.085 3.060 14.445 4.230 ;
        RECT  14.310 3.825 14.760 4.275 ;
        RECT  13.725 8.730 16.245 9.090 ;
        RECT  13.725 8.685 14.175 9.135 ;
        RECT  15.795 8.685 16.245 9.135 ;
    END
END drp_2

MACRO drp_1
    CLASS CORE ;
    FOREIGN drp_1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.440 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  17.370 6.975 18.810 7.335 ;
        RECT  18.450 4.095 18.810 7.335 ;
        RECT  16.830 4.095 18.810 4.455 ;
        RECT  17.865 2.160 18.225 4.455 ;
        RECT  17.370 6.975 17.730 9.270 ;
        END
    END q
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER metal1 ;
        RECT  3.060 4.680 3.420 5.040 ;
        END
    END ck
    PIN rb
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  14.175 7.155 14.445 7.425 ;
        RECT  7.740 7.155 8.010 7.425 ;
        RECT  1.485 7.155 1.755 7.425 ;
        LAYER metal2 ;
        RECT  14.085 7.065 14.535 7.515 ;
        RECT  1.395 7.110 14.535 7.470 ;
        RECT  7.650 7.065 8.100 7.515 ;
        RECT  1.395 7.065 1.845 7.515 ;
        LAYER metal1 ;
        RECT  14.085 7.065 14.535 7.515 ;
        RECT  7.650 7.065 8.100 7.515 ;
        RECT  1.395 7.065 1.845 7.515 ;
        END
    END rb
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 19.440 0.990 ;
        RECT  17.100 0.000 17.460 2.790 ;
        RECT  11.835 0.000 12.195 2.790 ;
        RECT  10.215 0.000 10.575 2.790 ;
        RECT  7.830 0.000 8.190 2.790 ;
        RECT  3.240 0.000 3.600 2.655 ;
        RECT  0.630 0.000 0.990 2.790 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 19.440 11.340 ;
        RECT  16.605 8.010 16.965 11.340 ;
        RECT  14.535 8.010 14.895 11.340 ;
        RECT  11.565 8.010 11.925 11.340 ;
        RECT  9.990 8.010 10.350 11.340 ;
        RECT  7.065 8.010 7.425 11.340 ;
        RECT  2.925 8.010 3.285 11.340 ;
        RECT  2.115 8.010 2.475 11.340 ;
        RECT  0.630 8.010 0.990 11.340 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  1.350 8.685 1.800 9.135 ;
        RECT  1.395 8.010 1.755 9.270 ;
        RECT  2.250 2.205 2.700 2.655 ;
        RECT  2.925 3.015 3.375 3.465 ;
        RECT  3.195 6.255 3.645 6.705 ;
        RECT  3.960 4.635 4.410 5.085 ;
        RECT  4.005 2.160 4.365 7.560 ;
        RECT  3.690 7.200 4.050 9.270 ;
        RECT  4.680 8.685 5.130 9.135 ;
        RECT  4.725 8.010 5.085 9.270 ;
        RECT  4.815 2.205 5.265 2.655 ;
        RECT  6.210 8.685 6.660 9.135 ;
        RECT  6.255 8.010 6.615 9.270 ;
        RECT  6.345 2.205 6.795 2.655 ;
        RECT  6.525 3.015 6.975 3.465 ;
        RECT  7.785 8.685 8.235 9.135 ;
        RECT  7.830 8.010 8.190 9.270 ;
        RECT  8.145 5.445 8.595 5.895 ;
        RECT  9.315 2.205 9.765 2.655 ;
        RECT  5.625 2.160 5.985 5.850 ;
        RECT  9.225 5.490 10.440 5.850 ;
        RECT  9.225 5.490 9.585 6.660 ;
        RECT  5.490 6.300 9.585 6.660 ;
        RECT  5.490 5.490 5.850 9.270 ;
        RECT  10.980 2.160 11.340 5.850 ;
        RECT  10.800 5.445 11.340 5.850 ;
        RECT  10.755 5.490 12.015 5.850 ;
        RECT  10.755 5.490 11.250 5.895 ;
        RECT  10.755 5.490 11.115 9.270 ;
        RECT  12.780 3.015 13.230 3.465 ;
        RECT  12.555 3.420 13.185 3.780 ;
        RECT  12.555 3.420 12.915 5.085 ;
        RECT  12.510 4.635 12.960 5.085 ;
        RECT  12.600 2.295 13.680 2.655 ;
        RECT  13.320 6.255 13.770 6.705 ;
        RECT  13.725 8.685 14.175 9.135 ;
        RECT  13.770 8.010 14.130 9.270 ;
        RECT  14.310 3.825 14.760 4.275 ;
        RECT  15.795 8.685 16.245 9.135 ;
        RECT  15.840 8.010 16.200 9.270 ;
        RECT  15.435 2.295 16.695 2.655 ;
        RECT  14.085 2.160 14.445 3.420 ;
        RECT  13.590 3.060 14.445 3.420 ;
        RECT  13.590 3.060 13.950 5.850 ;
        RECT  12.465 5.490 17.280 5.850 ;
        RECT  12.465 5.490 12.825 7.470 ;
        RECT  12.465 7.110 13.320 7.470 ;
        RECT  12.960 7.110 13.320 9.270 ;
        LAYER via ;
        RECT  1.440 8.775 1.710 9.045 ;
        RECT  2.340 2.295 2.610 2.565 ;
        RECT  3.015 3.105 3.285 3.375 ;
        RECT  3.285 6.345 3.555 6.615 ;
        RECT  4.050 4.725 4.320 4.995 ;
        RECT  4.770 8.775 5.040 9.045 ;
        RECT  4.905 2.295 5.175 2.565 ;
        RECT  6.300 8.775 6.570 9.045 ;
        RECT  6.435 2.295 6.705 2.565 ;
        RECT  6.615 3.105 6.885 3.375 ;
        RECT  7.875 8.775 8.145 9.045 ;
        RECT  8.235 5.535 8.505 5.805 ;
        RECT  9.405 2.295 9.675 2.565 ;
        RECT  10.890 5.535 11.160 5.805 ;
        RECT  12.600 4.725 12.870 4.995 ;
        RECT  12.870 3.105 13.140 3.375 ;
        RECT  13.410 6.345 13.680 6.615 ;
        RECT  13.815 8.775 14.085 9.045 ;
        RECT  14.400 3.915 14.670 4.185 ;
        RECT  15.885 8.775 16.155 9.045 ;
        LAYER metal2 ;
        RECT  1.350 8.730 5.130 9.090 ;
        RECT  1.350 8.685 1.800 9.135 ;
        RECT  4.680 8.685 5.130 9.135 ;
        RECT  2.250 2.250 5.265 2.610 ;
        RECT  2.250 2.205 2.700 2.655 ;
        RECT  4.815 2.205 5.265 2.655 ;
        RECT  2.925 3.060 6.975 3.420 ;
        RECT  2.925 3.015 3.375 3.465 ;
        RECT  6.525 3.015 6.975 3.465 ;
        RECT  6.210 8.730 8.235 9.090 ;
        RECT  6.210 8.685 6.660 9.135 ;
        RECT  7.785 8.685 8.235 9.135 ;
        RECT  6.345 2.250 9.765 2.610 ;
        RECT  6.345 2.205 6.795 2.655 ;
        RECT  9.315 2.205 9.765 2.655 ;
        RECT  8.145 5.490 11.250 5.850 ;
        RECT  8.145 5.445 8.595 5.895 ;
        RECT  10.800 5.445 11.250 5.895 ;
        RECT  3.960 4.680 12.960 5.040 ;
        RECT  3.960 4.635 4.410 5.085 ;
        RECT  12.510 4.635 12.960 5.085 ;
        RECT  3.195 6.300 13.770 6.660 ;
        RECT  3.195 6.255 3.645 6.705 ;
        RECT  13.320 6.255 13.770 6.705 ;
        RECT  12.780 3.060 14.445 3.420 ;
        RECT  12.780 3.015 13.230 3.465 ;
        RECT  14.085 3.060 14.445 4.230 ;
        RECT  14.310 3.825 14.760 4.275 ;
        RECT  13.725 8.730 16.245 9.090 ;
        RECT  13.725 8.685 14.175 9.135 ;
        RECT  15.795 8.685 16.245 9.135 ;
    END
END drp_1

MACRO dp_4
    CLASS CORE ;
    FOREIGN dp_4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.010 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER metal1 ;
        RECT  2.250 4.680 2.610 5.040 ;
        END
    END ck
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 3.870 0.990 4.230 ;
        END
    END ip
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  15.030 5.895 16.380 6.255 ;
        RECT  16.020 3.960 16.380 6.255 ;
        RECT  12.420 4.680 16.380 5.040 ;
        RECT  15.030 3.960 16.380 4.320 ;
        RECT  15.030 5.895 15.390 9.270 ;
        RECT  15.030 2.160 15.390 4.320 ;
        END
    END q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 17.010 11.340 ;
        RECT  15.795 6.750 16.155 11.340 ;
        RECT  14.265 6.750 14.625 11.340 ;
        RECT  12.600 8.010 12.960 11.340 ;
        RECT  9.765 8.010 10.125 11.340 ;
        RECT  8.190 8.010 8.550 11.340 ;
        RECT  6.030 8.010 6.390 11.340 ;
        RECT  2.250 8.010 2.610 11.340 ;
        RECT  0.630 8.010 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 17.010 0.990 ;
        RECT  15.840 0.000 16.200 3.420 ;
        RECT  14.220 0.000 14.580 3.420 ;
        RECT  13.410 0.000 13.770 2.790 ;
        RECT  9.765 0.000 10.125 2.790 ;
        RECT  8.190 0.000 8.550 2.790 ;
        RECT  6.300 0.000 6.660 2.700 ;
        RECT  2.250 0.000 2.610 2.700 ;
        RECT  0.630 0.000 0.990 2.790 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  1.350 8.685 1.800 9.135 ;
        RECT  1.395 8.010 1.755 9.270 ;
        RECT  1.350 2.205 1.800 2.655 ;
        RECT  1.935 3.015 2.385 3.465 ;
        RECT  2.610 6.255 3.060 6.705 ;
        RECT  3.015 2.160 3.375 3.420 ;
        RECT  3.015 3.060 3.870 3.420 ;
        RECT  3.465 4.635 3.915 5.085 ;
        RECT  3.510 3.060 3.870 7.650 ;
        RECT  3.060 7.290 3.870 7.650 ;
        RECT  3.060 7.290 3.420 9.270 ;
        RECT  3.825 2.205 4.275 2.655 ;
        RECT  3.915 8.685 4.365 9.135 ;
        RECT  3.960 8.010 4.320 9.270 ;
        RECT  5.355 2.205 5.805 2.655 ;
        RECT  5.805 5.445 6.255 5.895 ;
        RECT  5.850 3.015 6.300 3.465 ;
        RECT  6.975 2.205 7.425 2.655 ;
        RECT  4.635 2.160 4.995 5.670 ;
        RECT  7.650 5.490 8.775 5.850 ;
        RECT  7.650 5.490 8.010 6.840 ;
        RECT  4.725 6.480 8.010 6.840 ;
        RECT  4.725 5.220 5.085 9.270 ;
        RECT  8.955 2.160 9.315 3.465 ;
        RECT  9.090 5.490 10.305 5.850 ;
        RECT  9.090 5.445 9.540 5.895 ;
        RECT  9.135 3.105 9.495 7.650 ;
        RECT  8.955 7.290 9.315 9.270 ;
        RECT  10.710 3.015 11.160 3.465 ;
        RECT  10.755 3.015 11.115 5.085 ;
        RECT  10.710 4.635 11.160 5.085 ;
        RECT  10.485 2.295 11.565 2.655 ;
        RECT  11.520 6.255 11.970 6.705 ;
        RECT  12.645 3.015 13.095 3.465 ;
        RECT  12.690 3.015 13.050 4.275 ;
        RECT  12.375 3.915 13.050 4.275 ;
        RECT  11.970 2.160 12.330 3.420 ;
        RECT  11.565 3.060 12.330 3.420 ;
        RECT  11.565 3.060 11.925 5.850 ;
        RECT  10.710 5.490 14.760 5.850 ;
        RECT  10.710 5.490 11.070 7.650 ;
        RECT  10.710 7.290 11.475 7.650 ;
        RECT  11.115 7.290 11.475 9.270 ;
        LAYER via ;
        RECT  1.440 8.775 1.710 9.045 ;
        RECT  1.440 2.295 1.710 2.565 ;
        RECT  2.025 3.105 2.295 3.375 ;
        RECT  2.700 6.345 2.970 6.615 ;
        RECT  3.555 4.725 3.825 4.995 ;
        RECT  3.915 2.295 4.185 2.565 ;
        RECT  4.005 8.775 4.275 9.045 ;
        RECT  5.445 2.295 5.715 2.565 ;
        RECT  5.895 5.535 6.165 5.805 ;
        RECT  5.940 3.105 6.210 3.375 ;
        RECT  7.065 2.295 7.335 2.565 ;
        RECT  9.180 5.535 9.450 5.805 ;
        RECT  10.800 4.725 11.070 4.995 ;
        RECT  10.800 3.105 11.070 3.375 ;
        RECT  11.610 6.345 11.880 6.615 ;
        RECT  12.735 3.105 13.005 3.375 ;
        LAYER metal2 ;
        RECT  1.350 2.250 4.275 2.610 ;
        RECT  1.350 2.205 1.800 2.655 ;
        RECT  3.825 2.205 4.275 2.655 ;
        RECT  1.350 8.730 4.365 9.090 ;
        RECT  1.350 8.685 1.800 9.135 ;
        RECT  3.915 8.685 4.365 9.135 ;
        RECT  1.935 3.060 6.300 3.420 ;
        RECT  1.935 3.015 2.385 3.465 ;
        RECT  5.850 3.015 6.300 3.465 ;
        RECT  5.355 2.250 7.425 2.610 ;
        RECT  5.355 2.205 5.805 2.655 ;
        RECT  6.975 2.205 7.425 2.655 ;
        RECT  5.805 5.490 9.540 5.850 ;
        RECT  5.805 5.445 6.255 5.895 ;
        RECT  9.090 5.445 9.540 5.895 ;
        RECT  3.465 4.680 11.160 5.040 ;
        RECT  3.465 4.635 3.915 5.085 ;
        RECT  10.710 4.635 11.160 5.085 ;
        RECT  2.610 6.300 11.970 6.660 ;
        RECT  2.610 6.255 3.060 6.705 ;
        RECT  11.520 6.255 11.970 6.705 ;
        RECT  10.710 3.060 13.095 3.420 ;
        RECT  10.710 3.015 11.160 3.465 ;
        RECT  12.645 3.015 13.095 3.465 ;
    END
END dp_4

MACRO dp_2
    CLASS CORE ;
    FOREIGN dp_2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.200 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER metal1 ;
        RECT  2.250 4.680 2.610 5.040 ;
        END
    END ck
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.420 4.680 15.570 5.040 ;
        RECT  15.030 3.825 15.570 5.040 ;
        RECT  15.030 2.160 15.390 9.270 ;
        END
    END q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 16.200 0.990 ;
        RECT  14.220 0.000 14.580 3.420 ;
        RECT  13.410 0.000 13.770 2.790 ;
        RECT  9.765 0.000 10.125 2.790 ;
        RECT  8.190 0.000 8.550 2.790 ;
        RECT  6.300 0.000 6.660 2.700 ;
        RECT  2.250 0.000 2.610 2.700 ;
        RECT  0.630 0.000 0.990 2.790 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 16.200 11.340 ;
        RECT  14.265 6.750 14.625 11.340 ;
        RECT  12.600 8.010 12.960 11.340 ;
        RECT  9.765 8.010 10.125 11.340 ;
        RECT  8.190 8.010 8.550 11.340 ;
        RECT  6.030 8.010 6.390 11.340 ;
        RECT  2.250 8.010 2.610 11.340 ;
        RECT  0.630 8.010 0.990 11.340 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  1.350 8.685 1.800 9.135 ;
        RECT  1.395 8.010 1.755 9.270 ;
        RECT  1.350 2.205 1.800 2.655 ;
        RECT  1.935 3.015 2.385 3.465 ;
        RECT  2.610 6.255 3.060 6.705 ;
        RECT  3.015 2.160 3.375 3.465 ;
        RECT  3.015 3.105 3.870 3.465 ;
        RECT  3.465 4.635 3.915 5.085 ;
        RECT  3.510 3.105 3.870 7.650 ;
        RECT  3.060 7.290 3.870 7.650 ;
        RECT  3.060 7.290 3.420 9.270 ;
        RECT  3.825 2.205 4.275 2.655 ;
        RECT  3.915 8.685 4.365 9.135 ;
        RECT  3.960 8.010 4.320 9.270 ;
        RECT  5.355 2.205 5.805 2.655 ;
        RECT  5.805 5.445 6.255 5.895 ;
        RECT  5.850 3.015 6.300 3.465 ;
        RECT  6.975 2.205 7.425 2.655 ;
        RECT  4.635 2.160 4.995 5.670 ;
        RECT  7.650 5.490 8.775 5.850 ;
        RECT  7.650 5.490 8.010 6.840 ;
        RECT  4.725 6.480 8.010 6.840 ;
        RECT  4.725 5.220 5.085 9.270 ;
        RECT  8.955 2.160 9.315 3.465 ;
        RECT  9.090 5.490 10.305 5.850 ;
        RECT  9.090 5.445 9.540 5.895 ;
        RECT  9.135 3.105 9.495 7.650 ;
        RECT  8.955 7.290 9.315 9.270 ;
        RECT  10.710 3.015 11.160 3.465 ;
        RECT  10.755 3.015 11.115 5.085 ;
        RECT  10.710 4.635 11.160 5.085 ;
        RECT  10.485 2.295 11.565 2.655 ;
        RECT  11.520 6.255 11.970 6.705 ;
        RECT  12.330 3.825 12.780 4.275 ;
        RECT  11.970 2.160 12.330 3.465 ;
        RECT  11.565 3.105 12.330 3.465 ;
        RECT  11.565 3.105 11.925 5.850 ;
        RECT  10.710 5.490 14.760 5.850 ;
        RECT  10.710 5.490 11.070 7.650 ;
        RECT  10.710 7.290 11.475 7.650 ;
        RECT  11.115 7.290 11.475 9.270 ;
        LAYER via ;
        RECT  1.440 8.775 1.710 9.045 ;
        RECT  1.440 2.295 1.710 2.565 ;
        RECT  2.025 3.105 2.295 3.375 ;
        RECT  2.700 6.345 2.970 6.615 ;
        RECT  3.555 4.725 3.825 4.995 ;
        RECT  3.915 2.295 4.185 2.565 ;
        RECT  4.005 8.775 4.275 9.045 ;
        RECT  5.445 2.295 5.715 2.565 ;
        RECT  5.895 5.535 6.165 5.805 ;
        RECT  5.940 3.105 6.210 3.375 ;
        RECT  7.065 2.295 7.335 2.565 ;
        RECT  9.180 5.535 9.450 5.805 ;
        RECT  10.800 4.725 11.070 4.995 ;
        RECT  10.800 3.105 11.070 3.375 ;
        RECT  11.610 6.345 11.880 6.615 ;
        RECT  12.420 3.915 12.690 4.185 ;
        LAYER metal2 ;
        RECT  1.350 2.250 4.275 2.610 ;
        RECT  1.350 2.205 1.800 2.655 ;
        RECT  3.825 2.205 4.275 2.655 ;
        RECT  1.350 8.730 4.365 9.090 ;
        RECT  1.350 8.685 1.800 9.135 ;
        RECT  3.915 8.685 4.365 9.135 ;
        RECT  1.935 3.060 6.300 3.420 ;
        RECT  1.935 3.015 2.385 3.465 ;
        RECT  5.850 3.015 6.300 3.465 ;
        RECT  5.355 2.250 7.425 2.610 ;
        RECT  5.355 2.205 5.805 2.655 ;
        RECT  6.975 2.205 7.425 2.655 ;
        RECT  5.805 5.490 9.540 5.850 ;
        RECT  5.805 5.445 6.255 5.895 ;
        RECT  9.090 5.445 9.540 5.895 ;
        RECT  3.465 4.680 11.160 5.040 ;
        RECT  3.465 4.635 3.915 5.085 ;
        RECT  10.710 4.635 11.160 5.085 ;
        RECT  2.610 6.300 11.970 6.660 ;
        RECT  2.610 6.255 3.060 6.705 ;
        RECT  11.520 6.255 11.970 6.705 ;
        RECT  10.710 3.060 12.735 3.420 ;
        RECT  10.710 3.015 11.160 3.465 ;
        RECT  12.375 3.060 12.735 4.275 ;
        RECT  12.330 3.825 12.780 4.275 ;
    END
END dp_2

MACRO dp_1
    CLASS CORE ;
    FOREIGN dp_1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.390 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER metal1 ;
        RECT  2.250 4.680 2.610 5.040 ;
        END
    END ck
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.365 6.345 14.760 6.705 ;
        RECT  14.400 3.060 14.760 6.705 ;
        RECT  14.265 2.160 14.625 3.420 ;
        RECT  12.420 4.680 14.760 5.040 ;
        RECT  13.365 6.345 13.725 9.270 ;
        END
    END q
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 15.390 0.990 ;
        RECT  13.410 0.000 13.770 2.790 ;
        RECT  9.765 0.000 10.125 2.790 ;
        RECT  8.190 0.000 8.550 2.790 ;
        RECT  6.300 0.000 6.660 2.700 ;
        RECT  2.250 0.000 2.610 2.700 ;
        RECT  0.630 0.000 0.990 2.790 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 15.390 11.340 ;
        RECT  12.600 8.010 12.960 11.340 ;
        RECT  9.765 8.010 10.125 11.340 ;
        RECT  8.190 8.010 8.550 11.340 ;
        RECT  6.030 8.010 6.390 11.340 ;
        RECT  2.250 8.010 2.610 11.340 ;
        RECT  0.630 8.010 0.990 11.340 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  1.350 8.685 1.800 9.135 ;
        RECT  1.395 8.010 1.755 9.270 ;
        RECT  1.350 2.205 1.800 2.655 ;
        RECT  1.935 3.015 2.385 3.465 ;
        RECT  2.610 6.255 3.060 6.705 ;
        RECT  3.015 2.160 3.375 3.465 ;
        RECT  3.015 3.105 3.870 3.465 ;
        RECT  3.465 4.635 3.915 5.085 ;
        RECT  3.510 3.105 3.870 7.650 ;
        RECT  3.060 7.290 3.870 7.650 ;
        RECT  3.060 7.290 3.420 9.270 ;
        RECT  3.825 2.205 4.275 2.655 ;
        RECT  3.915 8.685 4.365 9.135 ;
        RECT  3.960 8.010 4.320 9.270 ;
        RECT  5.355 2.205 5.805 2.655 ;
        RECT  5.805 5.445 6.255 5.895 ;
        RECT  5.850 3.015 6.300 3.465 ;
        RECT  6.975 2.205 7.425 2.655 ;
        RECT  4.635 2.160 4.995 5.670 ;
        RECT  7.650 5.490 8.775 5.850 ;
        RECT  7.650 5.490 8.010 6.840 ;
        RECT  4.725 6.480 8.010 6.840 ;
        RECT  4.725 5.220 5.085 9.270 ;
        RECT  8.955 2.160 9.315 3.465 ;
        RECT  9.090 5.490 10.305 5.850 ;
        RECT  9.090 5.445 9.540 5.895 ;
        RECT  9.135 3.105 9.495 7.650 ;
        RECT  8.955 7.290 9.315 9.270 ;
        RECT  10.710 3.015 11.160 3.465 ;
        RECT  10.755 3.015 11.115 5.085 ;
        RECT  10.710 4.635 11.160 5.085 ;
        RECT  10.485 2.295 11.565 2.655 ;
        RECT  11.520 6.255 11.970 6.705 ;
        RECT  12.330 3.825 12.780 4.275 ;
        RECT  11.970 2.160 12.330 3.465 ;
        RECT  11.565 3.105 12.330 3.465 ;
        RECT  11.565 3.105 11.925 5.850 ;
        RECT  10.710 5.490 13.635 5.850 ;
        RECT  10.710 5.490 11.070 7.650 ;
        RECT  10.710 7.290 11.475 7.650 ;
        RECT  11.115 7.290 11.475 9.270 ;
        LAYER via ;
        RECT  1.440 8.775 1.710 9.045 ;
        RECT  1.440 2.295 1.710 2.565 ;
        RECT  2.025 3.105 2.295 3.375 ;
        RECT  2.700 6.345 2.970 6.615 ;
        RECT  3.555 4.725 3.825 4.995 ;
        RECT  3.915 2.295 4.185 2.565 ;
        RECT  4.005 8.775 4.275 9.045 ;
        RECT  5.445 2.295 5.715 2.565 ;
        RECT  5.895 5.535 6.165 5.805 ;
        RECT  5.940 3.105 6.210 3.375 ;
        RECT  7.065 2.295 7.335 2.565 ;
        RECT  9.180 5.535 9.450 5.805 ;
        RECT  10.800 4.725 11.070 4.995 ;
        RECT  10.800 3.105 11.070 3.375 ;
        RECT  11.610 6.345 11.880 6.615 ;
        RECT  12.420 3.915 12.690 4.185 ;
        LAYER metal2 ;
        RECT  1.350 2.250 4.275 2.610 ;
        RECT  1.350 2.205 1.800 2.655 ;
        RECT  3.825 2.205 4.275 2.655 ;
        RECT  1.350 8.730 4.365 9.090 ;
        RECT  1.350 8.685 1.800 9.135 ;
        RECT  3.915 8.685 4.365 9.135 ;
        RECT  1.935 3.060 6.300 3.420 ;
        RECT  1.935 3.015 2.385 3.465 ;
        RECT  5.850 3.015 6.300 3.465 ;
        RECT  5.355 2.250 7.425 2.610 ;
        RECT  5.355 2.205 5.805 2.655 ;
        RECT  6.975 2.205 7.425 2.655 ;
        RECT  5.805 5.490 9.540 5.850 ;
        RECT  5.805 5.445 6.255 5.895 ;
        RECT  9.090 5.445 9.540 5.895 ;
        RECT  3.465 4.680 11.160 5.040 ;
        RECT  3.465 4.635 3.915 5.085 ;
        RECT  10.710 4.635 11.160 5.085 ;
        RECT  2.610 6.300 11.970 6.660 ;
        RECT  2.610 6.255 3.060 6.705 ;
        RECT  11.520 6.255 11.970 6.705 ;
        RECT  10.710 3.060 12.735 3.420 ;
        RECT  10.710 3.015 11.160 3.465 ;
        RECT  12.375 3.060 12.735 4.275 ;
        RECT  12.330 3.825 12.780 4.275 ;
    END
END dp_1

MACRO dksp_1
    CLASS CORE ;
    FOREIGN dksp_1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 23.490 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN sb
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  3.060 3.870 3.420 4.230 ;
        END
    END sb
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip
    PIN qb
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  20.475 4.680 21.195 5.040 ;
        RECT  20.475 2.160 20.835 9.270 ;
        END
    END qb
    PIN ck
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER metal1 ;
        RECT  9.540 4.680 9.900 5.040 ;
        END
    END ck
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  22.005 4.680 22.860 5.040 ;
        RECT  22.005 2.160 22.365 9.270 ;
        END
    END q
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 23.490 11.340 ;
        RECT  21.240 6.750 21.600 11.340 ;
        RECT  19.755 6.750 20.115 11.340 ;
        RECT  18.270 8.010 18.630 11.340 ;
        RECT  16.785 8.010 17.145 11.340 ;
        RECT  11.520 8.010 11.880 11.340 ;
        RECT  10.035 8.010 10.395 11.340 ;
        RECT  8.460 8.010 8.820 11.340 ;
        RECT  6.975 8.010 7.335 11.340 ;
        RECT  3.600 8.010 3.960 11.340 ;
        RECT  2.115 8.010 2.475 11.340 ;
        RECT  0.630 8.010 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 23.490 0.990 ;
        RECT  21.240 0.000 21.600 3.420 ;
        RECT  19.755 0.000 20.115 3.420 ;
        RECT  18.270 0.000 18.630 2.790 ;
        RECT  16.785 0.000 17.145 2.790 ;
        RECT  11.520 0.000 11.880 2.790 ;
        RECT  10.035 0.000 10.395 2.790 ;
        RECT  8.460 0.000 8.820 2.790 ;
        RECT  6.975 0.000 7.335 2.790 ;
        RECT  2.160 0.000 2.520 2.790 ;
        RECT  0.630 0.000 0.990 2.790 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  1.395 6.615 1.980 6.975 ;
        RECT  1.395 2.160 1.755 9.270 ;
        RECT  3.645 2.160 4.725 2.520 ;
        RECT  4.365 2.160 4.725 3.150 ;
        RECT  3.645 2.160 4.005 3.600 ;
        RECT  3.690 3.240 4.050 5.850 ;
        RECT  2.880 5.490 4.725 5.850 ;
        RECT  2.880 5.490 3.240 9.270 ;
        RECT  4.365 5.490 4.725 9.270 ;
        RECT  4.320 3.825 4.770 4.275 ;
        RECT  5.130 6.255 5.580 6.705 ;
        RECT  5.175 2.160 5.535 9.270 ;
        RECT  5.850 7.065 6.300 7.515 ;
        RECT  5.895 2.160 6.255 9.270 ;
        RECT  6.525 5.445 6.975 5.895 ;
        RECT  6.525 3.825 6.975 4.275 ;
        RECT  6.885 6.255 7.335 6.705 ;
        RECT  7.740 4.680 8.370 5.040 ;
        RECT  7.695 6.255 8.145 6.705 ;
        RECT  7.740 2.160 8.100 9.270 ;
        RECT  9.225 2.160 9.585 4.410 ;
        RECT  8.730 4.050 9.585 4.410 ;
        RECT  8.730 4.050 9.090 5.670 ;
        RECT  8.730 5.310 9.585 5.670 ;
        RECT  9.180 7.065 9.630 7.515 ;
        RECT  9.225 5.310 9.585 9.270 ;
        RECT  10.755 3.015 11.205 3.465 ;
        RECT  10.800 4.680 11.880 5.040 ;
        RECT  10.755 5.445 11.205 5.895 ;
        RECT  10.755 7.065 11.205 7.515 ;
        RECT  10.800 2.160 11.160 9.270 ;
        RECT  12.240 3.825 12.690 4.275 ;
        RECT  12.285 2.160 12.645 9.270 ;
        RECT  13.095 7.065 13.545 7.515 ;
        RECT  13.770 3.825 14.220 4.275 ;
        RECT  13.905 2.160 14.265 3.150 ;
        RECT  13.140 2.790 14.265 3.150 ;
        RECT  13.140 2.790 13.500 5.850 ;
        RECT  13.140 5.490 14.265 5.850 ;
        RECT  13.860 6.255 14.310 6.705 ;
        RECT  13.905 5.490 14.265 9.270 ;
        RECT  14.670 4.635 15.615 5.085 ;
        RECT  14.670 2.160 15.030 9.270 ;
        RECT  15.390 3.825 15.840 4.275 ;
        RECT  15.435 2.160 15.795 3.150 ;
        RECT  15.435 2.790 16.470 3.150 ;
        RECT  15.975 5.445 16.470 5.895 ;
        RECT  16.110 2.790 16.470 5.895 ;
        RECT  15.435 5.535 16.470 5.895 ;
        RECT  15.435 5.535 15.795 9.270 ;
        RECT  16.785 4.635 17.235 5.085 ;
        RECT  17.550 3.555 18.765 3.915 ;
        RECT  17.550 2.160 17.910 9.270 ;
        RECT  18.990 5.445 19.440 5.895 ;
        RECT  19.035 2.160 19.395 9.270 ;
        RECT  21.195 5.445 21.645 5.895 ;
        LAYER via ;
        RECT  4.410 3.915 4.680 4.185 ;
        RECT  5.220 6.345 5.490 6.615 ;
        RECT  5.940 7.155 6.210 7.425 ;
        RECT  6.615 5.535 6.885 5.805 ;
        RECT  6.615 3.915 6.885 4.185 ;
        RECT  6.975 6.345 7.245 6.615 ;
        RECT  7.785 6.345 8.055 6.615 ;
        RECT  9.270 7.155 9.540 7.425 ;
        RECT  10.845 7.155 11.115 7.425 ;
        RECT  10.845 5.535 11.115 5.805 ;
        RECT  10.845 3.105 11.115 3.375 ;
        RECT  12.330 3.915 12.600 4.185 ;
        RECT  13.185 7.155 13.455 7.425 ;
        RECT  13.860 3.915 14.130 4.185 ;
        RECT  13.950 6.345 14.220 6.615 ;
        RECT  15.255 4.725 15.525 4.995 ;
        RECT  15.480 3.915 15.750 4.185 ;
        RECT  16.065 5.535 16.335 5.805 ;
        RECT  16.875 4.725 17.145 4.995 ;
        RECT  19.080 5.535 19.350 5.805 ;
        RECT  21.285 5.535 21.555 5.805 ;
        LAYER metal2 ;
        RECT  5.130 6.300 7.335 6.660 ;
        RECT  5.130 6.255 5.580 6.705 ;
        RECT  6.885 6.255 7.335 6.705 ;
        RECT  5.850 7.110 9.630 7.470 ;
        RECT  5.850 7.065 6.300 7.515 ;
        RECT  9.180 7.065 9.630 7.515 ;
        RECT  6.525 5.490 11.205 5.850 ;
        RECT  6.525 5.445 6.975 5.895 ;
        RECT  10.755 5.445 11.205 5.895 ;
        RECT  10.755 7.110 13.545 7.470 ;
        RECT  10.755 7.065 11.205 7.515 ;
        RECT  13.095 7.065 13.545 7.515 ;
        RECT  6.525 3.870 14.220 4.230 ;
        RECT  6.525 3.825 6.975 4.275 ;
        RECT  12.240 3.825 12.690 4.275 ;
        RECT  13.770 3.825 14.220 4.275 ;
        RECT  7.695 6.300 14.310 6.660 ;
        RECT  7.695 6.255 8.145 6.705 ;
        RECT  13.860 6.255 14.310 6.705 ;
        RECT  4.365 3.060 15.795 3.420 ;
        RECT  10.755 3.015 11.205 3.465 ;
        RECT  4.365 3.060 4.725 4.275 ;
        RECT  15.435 3.060 15.795 4.275 ;
        RECT  4.320 3.825 4.770 4.275 ;
        RECT  15.390 3.825 15.840 4.275 ;
        RECT  15.165 4.680 17.235 5.040 ;
        RECT  15.165 4.635 15.615 5.085 ;
        RECT  16.785 4.635 17.235 5.085 ;
        RECT  15.975 5.490 21.645 5.850 ;
        RECT  15.975 5.445 16.425 5.895 ;
        RECT  18.990 5.445 19.440 5.895 ;
        RECT  21.195 5.445 21.645 5.895 ;
    END
END dksp_1

MACRO cd_8
    CLASS CORE ;
    FOREIGN cd_8 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.100 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.850 6.120 7.470 6.480 ;
        RECT  7.110 3.780 7.470 6.480 ;
        RECT  5.850 3.780 7.470 4.140 ;
        RECT  5.850 6.120 6.210 9.270 ;
        RECT  5.850 2.160 6.210 4.140 ;
        END
    END op
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 8.100 0.990 ;
        RECT  6.570 0.000 6.930 3.420 ;
        RECT  5.085 0.000 5.445 3.420 ;
        RECT  3.600 0.000 3.960 3.420 ;
        RECT  2.115 0.000 2.475 3.420 ;
        RECT  0.630 0.000 0.990 3.420 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 8.100 11.340 ;
        RECT  6.570 6.750 6.930 11.340 ;
        RECT  5.085 6.750 5.445 11.340 ;
        RECT  3.600 6.750 3.960 11.340 ;
        RECT  2.115 6.750 2.475 11.340 ;
        RECT  0.630 6.750 0.990 11.340 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  1.395 5.490 2.970 5.850 ;
        RECT  1.395 2.160 1.755 9.270 ;
        RECT  2.880 2.160 3.240 4.140 ;
        RECT  2.880 3.780 3.690 4.140 ;
        RECT  3.330 5.490 4.455 5.850 ;
        RECT  3.330 3.780 3.690 6.480 ;
        RECT  2.880 6.120 3.690 6.480 ;
        RECT  2.880 6.120 3.240 9.270 ;
        RECT  4.365 2.160 4.725 4.140 ;
        RECT  4.365 3.780 5.175 4.140 ;
        RECT  4.815 5.490 5.940 5.850 ;
        RECT  4.815 3.780 5.175 6.480 ;
        RECT  4.365 6.120 5.175 6.480 ;
        RECT  4.365 6.120 4.725 9.270 ;
    END
END cd_8

MACRO cd_16
    CLASS CORE ;
    FOREIGN cd_16 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.580 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.600 6.120 13.950 6.480 ;
        RECT  13.590 3.780 13.950 6.480 ;
        RECT  12.600 3.780 13.950 4.140 ;
        RECT  12.600 6.120 12.960 9.270 ;
        RECT  12.600 2.160 12.960 4.140 ;
        END
    END op
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 14.580 11.340 ;
        RECT  13.320 6.750 13.680 11.340 ;
        RECT  11.835 6.750 12.195 11.340 ;
        RECT  10.350 6.750 10.710 11.340 ;
        RECT  8.865 6.750 9.225 11.340 ;
        RECT  7.380 6.750 7.740 11.340 ;
        RECT  6.570 6.750 6.930 11.340 ;
        RECT  5.085 6.750 5.445 11.340 ;
        RECT  3.600 6.750 3.960 11.340 ;
        RECT  2.115 6.750 2.475 11.340 ;
        RECT  0.630 6.750 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 14.580 0.990 ;
        RECT  13.320 0.000 13.680 3.420 ;
        RECT  11.835 0.000 12.195 3.420 ;
        RECT  10.350 0.000 10.710 3.420 ;
        RECT  8.865 0.000 9.225 3.420 ;
        RECT  7.380 0.000 7.740 3.420 ;
        RECT  6.570 0.000 6.930 3.420 ;
        RECT  5.085 0.000 5.445 3.420 ;
        RECT  3.600 0.000 3.960 3.420 ;
        RECT  2.115 0.000 2.475 3.420 ;
        RECT  0.630 0.000 0.990 3.420 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  1.395 5.490 2.970 5.850 ;
        RECT  1.395 2.160 1.755 9.270 ;
        RECT  2.880 2.160 3.240 4.140 ;
        RECT  2.880 3.780 3.690 4.140 ;
        RECT  3.330 5.490 4.455 5.850 ;
        RECT  3.330 3.780 3.690 6.480 ;
        RECT  2.880 6.120 3.690 6.480 ;
        RECT  2.880 6.120 3.240 9.270 ;
        RECT  4.365 2.160 4.725 4.140 ;
        RECT  4.365 3.780 5.175 4.140 ;
        RECT  4.815 5.490 5.940 5.850 ;
        RECT  4.815 3.780 5.175 6.480 ;
        RECT  4.365 6.120 5.175 6.480 ;
        RECT  4.365 6.120 4.725 9.270 ;
        RECT  5.850 2.160 6.210 4.140 ;
        RECT  5.850 3.780 6.660 4.140 ;
        RECT  6.300 5.490 8.235 5.850 ;
        RECT  6.300 3.780 6.660 6.480 ;
        RECT  5.850 6.120 6.660 6.480 ;
        RECT  5.850 6.120 6.210 9.270 ;
        RECT  8.145 2.160 8.505 4.140 ;
        RECT  8.145 3.780 8.955 4.140 ;
        RECT  8.595 5.490 9.720 5.850 ;
        RECT  8.595 3.780 8.955 6.480 ;
        RECT  8.145 6.120 8.955 6.480 ;
        RECT  8.145 6.120 8.505 9.270 ;
        RECT  9.630 2.160 9.990 4.140 ;
        RECT  9.630 3.780 10.440 4.140 ;
        RECT  10.080 5.490 11.205 5.850 ;
        RECT  10.080 3.780 10.440 6.480 ;
        RECT  9.630 6.120 10.440 6.480 ;
        RECT  9.630 6.120 9.990 9.270 ;
        RECT  11.115 2.160 11.475 4.140 ;
        RECT  11.115 3.780 11.925 4.140 ;
        RECT  11.565 5.490 12.690 5.850 ;
        RECT  11.565 3.780 11.925 6.480 ;
        RECT  11.115 6.120 11.925 6.480 ;
        RECT  11.115 6.120 11.475 9.270 ;
    END
END cd_16

MACRO cd_12
    CLASS CORE ;
    FOREIGN cd_12 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.530 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.775 6.120 9.900 6.480 ;
        RECT  9.540 3.780 9.900 6.480 ;
        RECT  8.775 3.780 9.900 4.140 ;
        RECT  8.775 6.120 9.135 9.270 ;
        RECT  8.775 2.160 9.135 4.140 ;
        END
    END op
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 10.530 0.990 ;
        RECT  9.495 0.000 9.855 3.420 ;
        RECT  8.055 0.000 8.415 3.420 ;
        RECT  6.570 0.000 6.930 3.420 ;
        RECT  5.085 0.000 5.445 3.420 ;
        RECT  3.600 0.000 3.960 3.420 ;
        RECT  2.115 0.000 2.475 3.420 ;
        RECT  0.630 0.000 0.990 3.420 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 10.530 11.340 ;
        RECT  9.495 6.750 9.855 11.340 ;
        RECT  8.055 6.750 8.415 11.340 ;
        RECT  6.570 6.750 6.930 11.340 ;
        RECT  5.085 6.750 5.445 11.340 ;
        RECT  3.600 6.750 3.960 11.340 ;
        RECT  2.115 6.750 2.475 11.340 ;
        RECT  0.630 6.750 0.990 11.340 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  1.395 5.490 2.970 5.850 ;
        RECT  1.395 2.160 1.755 9.270 ;
        RECT  2.880 2.160 3.240 4.140 ;
        RECT  2.880 3.780 3.690 4.140 ;
        RECT  3.330 5.490 4.455 5.850 ;
        RECT  3.330 3.780 3.690 6.480 ;
        RECT  2.880 6.120 3.690 6.480 ;
        RECT  2.880 6.120 3.240 9.270 ;
        RECT  4.365 2.160 4.725 4.140 ;
        RECT  4.365 3.780 5.175 4.140 ;
        RECT  4.815 5.490 5.940 5.850 ;
        RECT  4.815 3.780 5.175 6.480 ;
        RECT  4.365 6.120 5.175 6.480 ;
        RECT  4.365 6.120 4.725 9.270 ;
        RECT  5.850 2.160 6.210 4.140 ;
        RECT  5.850 3.780 6.660 4.140 ;
        RECT  6.300 5.490 7.425 5.850 ;
        RECT  6.300 3.780 6.660 6.480 ;
        RECT  5.850 6.120 6.660 6.480 ;
        RECT  5.850 6.120 6.210 9.270 ;
        RECT  7.335 2.160 7.695 4.140 ;
        RECT  7.335 3.780 8.145 4.140 ;
        RECT  7.785 5.490 8.910 5.850 ;
        RECT  7.785 3.780 8.145 6.480 ;
        RECT  7.335 6.120 8.145 6.480 ;
        RECT  7.335 6.120 7.695 9.270 ;
    END
END cd_12

MACRO bufzp_2
    CLASS CORE ;
    FOREIGN bufzp_2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.480 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.490 3.060 5.850 7.110 ;
        RECT  5.445 6.750 5.805 9.270 ;
        RECT  5.445 2.160 5.805 3.420 ;
        END
    END op
    PIN c
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER via ;
        RECT  4.725 5.535 4.995 5.805 ;
        RECT  2.295 5.535 2.565 5.805 ;
        LAYER metal2 ;
        RECT  4.635 5.445 5.085 5.895 ;
        RECT  2.205 5.490 5.085 5.850 ;
        RECT  2.205 5.445 2.655 5.895 ;
        LAYER metal1 ;
        RECT  4.635 5.445 5.085 5.895 ;
        RECT  2.205 5.445 2.655 5.895 ;
        RECT  2.250 4.680 2.610 5.895 ;
        END
    END c
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 6.480 11.340 ;
        RECT  3.870 6.750 4.230 11.340 ;
        RECT  2.250 8.010 2.610 11.340 ;
        RECT  0.630 8.010 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 6.480 0.990 ;
        RECT  3.870 0.000 4.230 3.420 ;
        RECT  2.250 0.000 2.610 2.790 ;
        RECT  0.630 0.000 0.990 2.790 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  1.395 3.825 1.845 4.275 ;
        RECT  1.395 2.160 1.755 9.270 ;
        RECT  3.015 4.635 3.465 5.085 ;
        RECT  3.015 2.160 3.375 9.270 ;
        RECT  3.825 3.825 4.275 4.275 ;
        RECT  4.635 4.635 5.085 5.085 ;
        LAYER via ;
        RECT  1.485 3.915 1.755 4.185 ;
        RECT  3.105 4.725 3.375 4.995 ;
        RECT  3.915 3.915 4.185 4.185 ;
        RECT  4.725 4.725 4.995 4.995 ;
        LAYER metal2 ;
        RECT  1.395 3.870 4.275 4.230 ;
        RECT  1.395 3.825 1.845 4.275 ;
        RECT  3.825 3.825 4.275 4.275 ;
        RECT  3.015 4.680 5.085 5.040 ;
        RECT  3.015 4.635 3.465 5.085 ;
        RECT  4.635 4.635 5.085 5.085 ;
    END
END bufzp_2

MACRO buf_4
    CLASS CORE ;
    FOREIGN buf_4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.860 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.835 5.490 4.230 5.850 ;
        RECT  3.870 3.870 4.230 5.850 ;
        RECT  2.835 3.870 4.230 4.230 ;
        RECT  2.835 5.490 3.195 9.270 ;
        RECT  2.835 2.160 3.195 4.230 ;
        END
    END op
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 4.860 11.340 ;
        RECT  3.555 6.750 3.915 11.340 ;
        RECT  2.115 6.750 2.475 11.340 ;
        RECT  0.630 6.750 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 4.860 0.990 ;
        RECT  3.555 0.000 3.915 3.420 ;
        RECT  2.115 0.000 2.475 3.420 ;
        RECT  0.630 0.000 0.990 3.420 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  1.395 4.680 2.925 5.040 ;
        RECT  1.395 2.160 1.755 9.270 ;
    END
END buf_4

MACRO buf_2
    CLASS CORE ;
    FOREIGN buf_2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.050 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.060 3.060 3.420 7.110 ;
        RECT  2.970 6.750 3.330 9.270 ;
        RECT  2.970 2.160 3.330 3.420 ;
        END
    END op
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 4.050 0.990 ;
        RECT  2.250 0.000 2.610 3.420 ;
        RECT  0.630 0.000 0.990 3.420 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 4.050 11.340 ;
        RECT  2.250 6.750 2.610 11.340 ;
        RECT  0.630 6.750 0.990 11.340 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  1.350 4.680 2.610 5.040 ;
        RECT  1.350 2.160 1.710 9.270 ;
    END
END buf_2

MACRO buf_1
    CLASS CORE ;
    FOREIGN buf_1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.050 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.970 3.870 3.420 4.230 ;
        RECT  2.970 2.160 3.330 9.270 ;
        END
    END op
    PIN ip
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 4.050 0.990 ;
        RECT  2.250 0.000 2.610 2.790 ;
        RECT  0.630 0.000 0.990 2.790 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 4.050 11.340 ;
        RECT  2.250 8.010 2.610 11.340 ;
        RECT  0.630 8.010 0.990 11.340 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  1.350 4.680 2.610 5.040 ;
        RECT  1.350 2.160 1.710 9.270 ;
    END
END buf_1

MACRO and4_4
    CLASS CORE ;
    FOREIGN and4_4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.480 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip1
    PIN ip3
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 4.680 2.610 5.040 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 5.490 2.610 5.850 ;
        END
    END ip2
    PIN ip4
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  3.060 3.870 3.420 4.230 ;
        END
    END ip4
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.680 5.490 5.850 5.850 ;
        RECT  5.490 3.870 5.850 5.850 ;
        RECT  4.680 3.870 5.850 4.230 ;
        RECT  4.680 5.490 5.040 9.270 ;
        RECT  4.680 2.160 5.040 4.230 ;
        END
    END op
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 6.480 11.340 ;
        RECT  5.490 6.750 5.850 11.340 ;
        RECT  3.870 6.750 4.230 11.340 ;
        RECT  2.250 7.470 2.610 11.340 ;
        RECT  0.630 6.750 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 6.480 0.990 ;
        RECT  5.490 0.000 5.850 3.420 ;
        RECT  3.870 0.000 4.230 3.420 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  0.630 2.160 0.990 5.085 ;
        RECT  0.630 4.680 1.800 5.040 ;
        RECT  0.630 4.635 1.080 5.085 ;
        RECT  1.440 6.300 3.420 6.660 ;
        RECT  1.440 4.680 1.800 9.270 ;
        RECT  3.060 6.300 3.420 9.270 ;
        RECT  4.230 4.635 4.680 5.085 ;
        LAYER via ;
        RECT  0.720 4.725 0.990 4.995 ;
        RECT  4.320 4.725 4.590 4.995 ;
        LAYER metal2 ;
        RECT  0.630 4.680 4.680 5.040 ;
        RECT  0.630 4.635 1.080 5.085 ;
        RECT  4.230 4.635 4.680 5.085 ;
    END
END and4_4

MACRO and4_2
    CLASS CORE ;
    FOREIGN and4_2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 5.490 2.610 5.850 ;
        END
    END ip2
    PIN ip4
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  3.060 3.870 3.420 4.230 ;
        END
    END ip4
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.680 2.160 5.040 9.270 ;
        END
    END op
    PIN ip3
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 4.680 2.610 5.040 ;
        END
    END ip3
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip1
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 5.670 11.340 ;
        RECT  3.870 6.750 4.230 11.340 ;
        RECT  2.250 7.290 2.610 11.340 ;
        RECT  0.630 6.750 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 5.670 0.990 ;
        RECT  3.870 0.000 4.230 3.420 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  0.630 2.160 0.990 5.085 ;
        RECT  0.630 4.680 1.800 5.040 ;
        RECT  0.630 4.635 1.080 5.085 ;
        RECT  1.440 6.300 3.420 6.660 ;
        RECT  1.440 4.680 1.800 9.270 ;
        RECT  3.060 6.300 3.420 9.270 ;
        RECT  3.960 4.635 4.410 5.085 ;
        LAYER via ;
        RECT  0.720 4.725 0.990 4.995 ;
        RECT  4.050 4.725 4.320 4.995 ;
        LAYER metal2 ;
        RECT  0.630 4.680 4.410 5.040 ;
        RECT  0.630 4.635 1.080 5.085 ;
        RECT  3.960 4.635 4.410 5.085 ;
    END
END and4_2

MACRO and4_1
    CLASS CORE ;
    FOREIGN and4_1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 6.300 0.990 6.660 ;
        END
    END ip1
    PIN ip3
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 5.490 2.610 5.850 ;
        END
    END ip3
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 3.870 1.800 4.230 ;
        END
    END ip2
    PIN ip4
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  3.060 3.060 3.420 3.420 ;
        END
    END ip4
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.680 2.160 5.040 9.270 ;
        END
    END op
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 5.670 11.340 ;
        RECT  3.870 7.920 4.230 11.340 ;
        RECT  2.250 7.920 2.610 11.340 ;
        RECT  0.630 7.920 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 5.670 0.990 ;
        RECT  3.870 0.000 4.230 2.790 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  0.630 2.160 0.990 5.040 ;
        RECT  0.630 4.680 4.230 5.040 ;
        RECT  1.440 7.110 3.420 7.470 ;
        RECT  1.440 4.680 1.800 9.270 ;
        RECT  3.060 7.110 3.420 9.270 ;
    END
END and4_1

MACRO and3_4
    CLASS CORE ;
    FOREIGN and3_4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.670 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 4.680 1.800 5.040 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip1
    PIN ip3
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  3.060 5.490 3.420 5.850 ;
        END
    END ip3
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.870 3.870 4.230 5.850 ;
        RECT  3.690 5.490 4.050 9.270 ;
        RECT  3.645 2.160 4.005 4.230 ;
        END
    END op
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 5.670 11.340 ;
        RECT  4.500 6.750 4.860 11.340 ;
        RECT  2.925 6.750 3.285 11.340 ;
        RECT  1.395 6.750 1.755 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 5.670 0.990 ;
        RECT  4.500 0.000 4.860 3.420 ;
        RECT  2.835 0.000 3.195 3.420 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  0.630 2.160 0.990 4.230 ;
        RECT  0.630 3.870 2.610 4.230 ;
        RECT  2.205 4.635 2.655 5.085 ;
        RECT  2.250 3.870 2.610 6.480 ;
        RECT  0.630 6.120 2.610 6.480 ;
        RECT  0.630 6.120 0.990 9.270 ;
        RECT  2.160 6.120 2.520 9.270 ;
        RECT  3.015 4.635 3.465 5.085 ;
        LAYER via ;
        RECT  2.295 4.725 2.565 4.995 ;
        RECT  3.105 4.725 3.375 4.995 ;
        LAYER metal2 ;
        RECT  2.205 4.680 3.465 5.040 ;
        RECT  2.205 4.635 2.655 5.085 ;
        RECT  3.015 4.635 3.465 5.085 ;
    END
END and3_4

MACRO and3_2
    CLASS CORE ;
    FOREIGN and3_2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.860 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.870 2.160 4.230 9.270 ;
        RECT  3.780 3.915 4.230 4.185 ;
        END
    END op
    PIN ip3
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  3.060 4.680 3.420 5.040 ;
        END
    END ip3
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip1
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 4.680 1.800 5.040 ;
        END
    END ip2
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 4.860 0.990 ;
        RECT  3.060 0.000 3.420 3.420 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 4.860 11.340 ;
        RECT  3.060 6.750 3.420 11.340 ;
        RECT  1.440 6.750 1.800 11.340 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  0.630 2.160 0.990 4.230 ;
        RECT  0.630 3.870 2.610 4.230 ;
        RECT  2.250 5.490 3.420 5.850 ;
        RECT  0.630 6.120 2.610 6.480 ;
        RECT  0.630 6.120 0.990 9.270 ;
        RECT  2.250 3.870 2.610 9.270 ;
    END
END and3_2

MACRO and3_1
    CLASS CORE ;
    FOREIGN and3_1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.860 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.870 2.160 4.230 9.270 ;
        END
    END op
    PIN ip3
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 6.390 2.610 6.750 ;
        END
    END ip3
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip1
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 3.870 1.800 4.230 ;
        END
    END ip2
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 4.860 0.990 ;
        RECT  3.060 0.000 3.420 2.790 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 4.860 11.340 ;
        RECT  3.060 8.010 3.420 11.340 ;
        RECT  1.440 8.010 1.800 11.340 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  0.630 2.160 0.990 5.040 ;
        RECT  0.630 4.680 3.420 5.040 ;
        RECT  1.440 4.680 1.800 7.470 ;
        RECT  0.630 7.110 2.610 7.470 ;
        RECT  0.630 7.110 0.990 9.270 ;
        RECT  2.250 7.110 2.610 9.270 ;
    END
END and3_1

MACRO and2_4
    CLASS CORE ;
    FOREIGN and2_4 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.860 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 4.680 1.800 5.040 ;
        END
    END ip2
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip1
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.060 2.160 3.420 9.270 ;
        END
    END op
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 4.860 11.340 ;
        RECT  3.870 6.750 4.230 11.340 ;
        RECT  2.250 6.750 2.610 11.340 ;
        RECT  0.630 6.750 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 4.860 0.990 ;
        RECT  3.870 0.000 4.230 3.420 ;
        RECT  2.250 0.000 2.610 3.420 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  0.630 2.160 0.990 4.230 ;
        RECT  0.630 3.870 2.610 4.230 ;
        RECT  2.250 3.870 2.610 5.850 ;
        RECT  1.440 5.490 2.610 5.850 ;
        RECT  1.440 5.490 1.800 9.270 ;
    END
END and2_4

MACRO and2_2
    CLASS CORE ;
    FOREIGN and2_2 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.050 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.060 2.160 3.420 9.270 ;
        END
    END op
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip1
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 4.680 1.800 5.040 ;
        END
    END ip2
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 4.050 0.990 ;
        RECT  2.250 0.000 2.610 3.420 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 4.050 11.340 ;
        RECT  2.250 6.750 2.610 11.340 ;
        RECT  0.630 6.750 0.990 11.340 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  0.630 2.160 0.990 4.230 ;
        RECT  0.630 3.870 2.610 4.230 ;
        RECT  2.250 3.870 2.610 5.850 ;
        RECT  1.440 5.490 2.610 5.850 ;
        RECT  1.440 5.490 1.800 9.270 ;
    END
END and2_2

MACRO and2_1
    CLASS CORE ;
    FOREIGN and2_1 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.050 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.060 2.160 3.420 9.270 ;
        END
    END op
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip1
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 4.680 1.800 5.040 ;
        END
    END ip2
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 4.050 0.990 ;
        RECT  2.250 0.000 2.610 2.790 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 4.050 11.340 ;
        RECT  2.250 8.010 2.610 11.340 ;
        RECT  0.630 8.010 0.990 11.340 ;
        END
    END vdd!
    OBS
        LAYER metal1 ;
        RECT  0.630 2.160 0.990 4.230 ;
        RECT  0.630 3.870 2.610 4.230 ;
        RECT  2.250 3.870 2.610 5.850 ;
        RECT  1.440 5.490 2.610 5.850 ;
        RECT  1.440 5.490 1.800 9.270 ;
    END
END and2_1

MACRO aborc
    CLASS CORE ;
    FOREIGN aborc 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.480 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 4.680 1.800 5.040 ;
        END
    END ip2
    PIN ip3
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 3.870 2.610 4.230 ;
        END
    END ip3
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip1
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.490 3.060 5.850 7.290 ;
        RECT  5.130 6.930 5.490 9.270 ;
        RECT  5.130 2.160 5.490 3.420 ;
        END
    END op
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 6.480 11.340 ;
        RECT  4.410 8.010 4.770 11.340 ;
        RECT  2.070 8.010 2.430 11.340 ;
        RECT  0.630 8.010 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 6.480 0.990 ;
        RECT  4.410 0.000 4.770 2.790 ;
        RECT  1.890 0.000 2.250 2.790 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  1.350 6.930 3.240 7.290 ;
        RECT  1.350 6.930 1.710 9.270 ;
        RECT  2.880 6.930 3.240 9.270 ;
        RECT  0.630 2.160 0.990 3.555 ;
        RECT  2.610 2.160 2.970 3.555 ;
        RECT  0.630 3.195 4.230 3.555 ;
        RECT  3.870 3.195 4.230 7.290 ;
        RECT  3.600 6.930 3.960 9.270 ;
    END
END aborc

MACRO abnorc
    CLASS CORE ;
    FOREIGN abnorc 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.860 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  1.440 4.680 1.800 5.040 ;
        END
    END ip2
    PIN ip3
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 3.870 2.610 4.230 ;
        END
    END ip3
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 5.490 0.990 5.850 ;
        END
    END ip1
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.870 3.195 4.230 7.290 ;
        RECT  3.600 6.930 3.960 9.270 ;
        RECT  0.630 3.195 4.230 3.555 ;
        RECT  2.610 2.160 2.970 3.555 ;
        RECT  0.630 2.160 0.990 3.555 ;
        END
    END op
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 4.860 11.340 ;
        RECT  2.070 8.010 2.430 11.340 ;
        RECT  0.630 8.010 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 4.860 0.990 ;
        RECT  1.890 0.000 2.250 2.790 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  1.350 6.930 3.240 7.290 ;
        RECT  1.350 6.930 1.710 9.270 ;
        RECT  2.880 6.930 3.240 9.270 ;
    END
END abnorc

MACRO ab_or_c_or_d
    CLASS CORE ;
    FOREIGN ab_or_c_or_d 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.290 BY 11.340 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN ip1
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  0.630 3.870 0.990 4.230 ;
        END
    END ip1
    PIN ip2
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  2.250 4.680 2.610 5.040 ;
        END
    END ip2
    PIN ip3
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  3.060 5.490 3.420 5.850 ;
        RECT  3.060 5.490 3.330 5.895 ;
        END
    END ip3
    PIN ip4
        DIRECTION INPUT ;
        USE ANALOG ;
        PORT
        LAYER metal1 ;
        RECT  4.680 3.870 5.040 4.230 ;
        END
    END ip4
    PIN op
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.300 2.160 6.660 9.270 ;
        END
    END op
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 10.350 7.290 11.340 ;
        RECT  5.490 8.010 5.850 11.340 ;
        RECT  2.250 8.010 2.610 11.340 ;
        RECT  0.630 8.010 0.990 11.340 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 0.000 7.290 0.990 ;
        RECT  5.490 0.000 5.850 2.790 ;
        RECT  4.680 0.000 5.040 2.790 ;
        RECT  3.060 0.000 3.420 2.790 ;
        RECT  0.630 0.000 0.990 2.790 ;
        END
    END gnd!
    OBS
        LAYER metal1 ;
        RECT  1.440 7.110 3.420 7.470 ;
        RECT  1.440 7.110 1.800 9.270 ;
        RECT  3.060 7.110 3.420 9.270 ;
        RECT  2.250 2.160 2.610 3.420 ;
        RECT  2.250 3.060 4.230 3.420 ;
        RECT  3.870 2.160 4.230 5.850 ;
        RECT  3.870 5.490 5.850 5.850 ;
        RECT  4.680 5.490 5.040 9.270 ;
    END
END ab_or_c_or_d

END LIBRARY
