
module vscale_alu ( op, in1, in2, out );
  input [3:0] op;
  input [31:0] in1;
  input [31:0] in2;
  output [31:0] out;
  wire   N316, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132;
  assign N316 = in1[31];

  inv_1 U831 ( .ip(op[1]), .op(n1771) );
  inv_1 U832 ( .ip(op[0]), .op(n1748) );
  inv_1 U833 ( .ip(op[3]), .op(n815) );
  nand2_1 U834 ( .ip1(n815), .ip2(op[2]), .op(n1176) );
  inv_1 U835 ( .ip(n1176), .op(n797) );
  nand3_1 U836 ( .ip1(n1771), .ip2(n1748), .ip3(n797), .op(n1985) );
  inv_1 U837 ( .ip(n1985), .op(n2096) );
  inv_1 U838 ( .ip(in1[30]), .op(n799) );
  nand2_1 U839 ( .ip1(in2[30]), .ip2(n799), .op(n1599) );
  nor2_1 U840 ( .ip1(in2[30]), .ip2(n799), .op(n1689) );
  inv_1 U841 ( .ip(n1689), .op(n1539) );
  nand2_1 U842 ( .ip1(n1599), .ip2(n1539), .op(n1715) );
  nor2_1 U843 ( .ip1(in2[30]), .ip2(in1[30]), .op(n798) );
  nor2_1 U844 ( .ip1(n1176), .ip2(n1771), .op(n2092) );
  inv_1 U845 ( .ip(n2092), .op(n1989) );
  nor2_1 U846 ( .ip1(op[0]), .ip2(n1989), .op(n2099) );
  inv_1 U847 ( .ip(n2099), .op(n2046) );
  nor2_1 U848 ( .ip1(n798), .ip2(n2046), .op(n802) );
  inv_1 U849 ( .ip(in2[30]), .op(n800) );
  nor3_1 U850 ( .ip1(n1989), .ip2(n800), .ip3(n799), .op(n801) );
  not_ab_or_c_or_d U851 ( .ip1(n2096), .ip2(n1715), .ip3(n802), .ip4(n801), 
        .op(n818) );
  inv_1 U852 ( .ip(op[2]), .op(n1696) );
  nand3_1 U853 ( .ip1(op[1]), .ip2(op[3]), .ip3(n1696), .op(n825) );
  inv_1 U854 ( .ip(n825), .op(n803) );
  nand2_1 U855 ( .ip1(op[0]), .ip2(n803), .op(n1198) );
  inv_1 U856 ( .ip(in2[4]), .op(n2100) );
  nor2_1 U857 ( .ip1(n1198), .ip2(n2100), .op(n1874) );
  nand2_1 U858 ( .ip1(n1874), .ip2(N316), .op(n2001) );
  nor2_1 U859 ( .ip1(in2[3]), .ip2(n1149), .op(n2022) );
  inv_1 U860 ( .ip(in1[7]), .op(n1376) );
  inv_1 U861 ( .ip(in2[0]), .op(n1772) );
  nor2_1 U862 ( .ip1(n1058), .ip2(n1772), .op(n1486) );
  inv_1 U863 ( .ip(n1486), .op(n1783) );
  nor2_1 U864 ( .ip1(n1376), .ip2(n1783), .op(n1441) );
  inv_1 U865 ( .ip(in1[9]), .op(n1389) );
  nand2_1 U866 ( .ip1(in2[0]), .ip2(n1058), .op(n2007) );
  nor2_1 U867 ( .ip1(n1389), .ip2(n2007), .op(n1363) );
  nand2_1 U868 ( .ip1(in2[1]), .ip2(n1772), .op(n2102) );
  inv_1 U869 ( .ip(n2102), .op(n1508) );
  nand2_1 U870 ( .ip1(in1[8]), .ip2(n1508), .op(n1417) );
  inv_1 U871 ( .ip(n1417), .op(n804) );
  inv_1 U872 ( .ip(in1[10]), .op(n1391) );
  nor2_1 U873 ( .ip1(in2[1]), .ip2(in2[0]), .op(n2048) );
  inv_1 U874 ( .ip(n2048), .op(n1782) );
  nor2_1 U875 ( .ip1(n1391), .ip2(n1782), .op(n1304) );
  or4_1 U876 ( .ip1(n1441), .ip2(n1363), .ip3(n804), .ip4(n1304), .op(n1906)
         );
  inv_1 U877 ( .ip(in1[5]), .op(n1857) );
  nor2_1 U878 ( .ip1(n1857), .ip2(n2007), .op(n1442) );
  nand2_1 U879 ( .ip1(in1[6]), .ip2(n2048), .op(n1418) );
  nand2_1 U880 ( .ip1(in1[3]), .ip2(n1486), .op(n805) );
  nand2_1 U881 ( .ip1(n1418), .ip2(n805), .op(n806) );
  not_ab_or_c_or_d U882 ( .ip1(n1508), .ip2(in1[4]), .ip3(n1442), .ip4(n806), 
        .op(n1904) );
  inv_1 U883 ( .ip(n2007), .op(n2106) );
  inv_1 U884 ( .ip(in1[2]), .op(n1472) );
  nor2_1 U885 ( .ip1(n1472), .ip2(n1782), .op(n808) );
  inv_1 U886 ( .ip(in1[0]), .op(n1770) );
  nor2_1 U887 ( .ip1(n1770), .ip2(n2102), .op(n807) );
  not_ab_or_c_or_d U888 ( .ip1(in1[1]), .ip2(n2106), .ip3(n808), .ip4(n807), 
        .op(n1927) );
  mux2_1 U889 ( .ip1(n1904), .ip2(n1927), .s(in2[2]), .op(n1406) );
  nor2_1 U890 ( .ip1(n1131), .ip2(n1406), .op(n814) );
  inv_1 U891 ( .ip(in1[12]), .op(n1661) );
  nand2_1 U892 ( .ip1(n1508), .ip2(n1661), .op(n812) );
  inv_1 U893 ( .ip(in1[14]), .op(n1882) );
  nand2_1 U894 ( .ip1(n2048), .ip2(n1882), .op(n811) );
  inv_1 U895 ( .ip(in1[11]), .op(n1359) );
  nand2_1 U896 ( .ip1(n1486), .ip2(n1359), .op(n810) );
  inv_1 U897 ( .ip(in1[13]), .op(n1554) );
  nand2_1 U898 ( .ip1(n2106), .ip2(n1554), .op(n809) );
  nand4_1 U899 ( .ip1(n812), .ip2(n811), .ip3(n810), .ip4(n809), .op(n989) );
  inv_1 U900 ( .ip(n1149), .op(n1509) );
  nor2_1 U901 ( .ip1(in2[3]), .ip2(n1509), .op(n2014) );
  inv_1 U902 ( .ip(n2014), .op(n2024) );
  nor2_1 U903 ( .ip1(n989), .ip2(n2024), .op(n813) );
  not_ab_or_c_or_d U904 ( .ip1(n2022), .ip2(n1906), .ip3(n814), .ip4(n813), 
        .op(n1886) );
  nand3_1 U905 ( .ip1(n1696), .ip2(n1771), .ip3(n815), .op(n826) );
  nor2_1 U906 ( .ip1(n826), .ip2(n1748), .op(n2124) );
  nand2_1 U907 ( .ip1(n2124), .ip2(in2[4]), .op(n2041) );
  or2_1 U908 ( .ip1(n1886), .ip2(n2041), .op(n817) );
  inv_1 U909 ( .ip(N316), .op(n2093) );
  nor2_1 U910 ( .ip1(n1198), .ip2(n2093), .op(n903) );
  nand2_1 U911 ( .ip1(n903), .ip2(n2024), .op(n816) );
  and4_1 U912 ( .ip1(n818), .ip2(n2001), .ip3(n817), .ip4(n816), .op(n855) );
  nor2_1 U913 ( .ip1(in2[4]), .ip2(n1198), .op(n1922) );
  nand2_1 U914 ( .ip1(N316), .ip2(in2[1]), .op(n886) );
  inv_1 U915 ( .ip(n886), .op(n820) );
  nor2_1 U916 ( .ip1(in1[30]), .ip2(in2[0]), .op(n819) );
  not_ab_or_c_or_d U917 ( .ip1(in2[0]), .ip2(n2093), .ip3(in2[1]), .ip4(n819), 
        .op(n1875) );
  nor2_1 U918 ( .ip1(n820), .ip2(n1875), .op(n984) );
  inv_1 U919 ( .ip(n984), .op(n1873) );
  nand2_1 U920 ( .ip1(n1922), .ip2(n1873), .op(n823) );
  nor3_1 U921 ( .ip1(op[1]), .ip2(n1748), .ip3(n1176), .op(n1214) );
  inv_1 U922 ( .ip(n1214), .op(n821) );
  nor2_1 U923 ( .ip1(in2[4]), .ip2(n821), .op(n2098) );
  nand2_1 U924 ( .ip1(n1875), .ip2(n2098), .op(n822) );
  nand2_1 U925 ( .ip1(n823), .ip2(n822), .op(n824) );
  nand2_1 U926 ( .ip1(n2014), .ip2(n824), .op(n854) );
  nor2_1 U927 ( .ip1(op[0]), .ip2(n825), .op(n1801) );
  xor2_1 U928 ( .ip1(n1801), .ip2(in2[30]), .op(n2088) );
  xor2_1 U929 ( .ip1(n1801), .ip2(in2[29]), .op(n2080) );
  xor2_1 U930 ( .ip1(n1801), .ip2(in2[28]), .op(n2039) );
  xor2_1 U931 ( .ip1(n1801), .ip2(in2[27]), .op(n1967) );
  xor2_1 U932 ( .ip1(n1801), .ip2(in2[26]), .op(n862) );
  xor2_1 U933 ( .ip1(n1801), .ip2(in2[25]), .op(n927) );
  xor2_1 U934 ( .ip1(n1801), .ip2(in2[24]), .op(n1934) );
  xor2_1 U935 ( .ip1(n1801), .ip2(in2[23]), .op(n963) );
  xor2_1 U936 ( .ip1(n1801), .ip2(in2[22]), .op(n996) );
  xor2_1 U937 ( .ip1(n1801), .ip2(in2[21]), .op(n1026) );
  xor2_1 U938 ( .ip1(n1801), .ip2(in2[20]), .op(n1040) );
  xor2_1 U939 ( .ip1(n1801), .ip2(in2[19]), .op(n1097) );
  xor2_1 U940 ( .ip1(n1801), .ip2(in2[18]), .op(n1925) );
  xor2_1 U941 ( .ip1(n1801), .ip2(in2[17]), .op(n1123) );
  buf_1 U942 ( .ip(n1801), .op(n2085) );
  xor2_1 U943 ( .ip1(n2085), .ip2(in2[16]), .op(n1148) );
  xor2_1 U944 ( .ip1(n2085), .ip2(in2[15]), .op(n1185) );
  xor2_1 U945 ( .ip1(n2085), .ip2(in2[14]), .op(n1895) );
  xor2_1 U946 ( .ip1(n2085), .ip2(in2[13]), .op(n1224) );
  xor2_1 U947 ( .ip1(n2085), .ip2(in2[12]), .op(n1250) );
  xor2_1 U948 ( .ip1(n2085), .ip2(in2[11]), .op(n1273) );
  xor2_1 U949 ( .ip1(n2085), .ip2(in2[10]), .op(n1294) );
  xor2_1 U950 ( .ip1(n2085), .ip2(in2[9]), .op(n1342) );
  xor2_1 U951 ( .ip1(n2085), .ip2(in2[8]), .op(n1357) );
  xor2_1 U952 ( .ip1(n2085), .ip2(in2[7]), .op(n1383) );
  xor2_1 U953 ( .ip1(n2085), .ip2(in2[6]), .op(n1426) );
  xor2_1 U954 ( .ip1(n2085), .ip2(in2[5]), .op(n1863) );
  xor2_1 U955 ( .ip1(n2085), .ip2(in2[4]), .op(n1456) );
  xor2_1 U956 ( .ip1(n2085), .ip2(in2[3]), .op(n1827) );
  xor2_1 U957 ( .ip1(n2085), .ip2(n1509), .op(n1464) );
  xor2_1 U958 ( .ip1(n2085), .ip2(in2[1]), .op(n1531) );
  xor2_1 U959 ( .ip1(n2085), .ip2(in2[0]), .op(n1800) );
  nor2_1 U960 ( .ip1(op[0]), .ip2(n826), .op(n827) );
  or2_1 U961 ( .ip1(n1801), .ip2(n827), .op(n2131) );
  nand2_1 U962 ( .ip1(n828), .ip2(n2131), .op(n853) );
  nand2_1 U963 ( .ip1(n2124), .ip2(n2100), .op(n1907) );
  inv_1 U964 ( .ip(n1907), .op(n2037) );
  inv_1 U965 ( .ip(in1[16]), .op(n1543) );
  inv_1 U966 ( .ip(in1[15]), .op(n1580) );
  mux2_1 U967 ( .ip1(n1543), .ip2(n1580), .s(in2[0]), .op(n1044) );
  nand2_1 U968 ( .ip1(in2[1]), .ip2(n1044), .op(n831) );
  or2_1 U969 ( .ip1(in1[18]), .ip2(in2[1]), .op(n829) );
  nand2_1 U970 ( .ip1(n829), .ip2(n2007), .op(n1297) );
  nand2_1 U971 ( .ip1(in2[0]), .ip2(in1[17]), .op(n1153) );
  nand2_1 U972 ( .ip1(n1297), .ip2(n1153), .op(n830) );
  nand2_1 U973 ( .ip1(n831), .ip2(n830), .op(n987) );
  nand2_1 U974 ( .ip1(in2[3]), .ip2(n1509), .op(n2003) );
  inv_1 U975 ( .ip(n2003), .op(n1946) );
  nand2_1 U976 ( .ip1(in1[27]), .ip2(in2[0]), .op(n2009) );
  inv_1 U977 ( .ip(in1[29]), .op(n2103) );
  nor2_1 U978 ( .ip1(n1772), .ip2(n2103), .op(n1064) );
  not_ab_or_c_or_d U979 ( .ip1(in1[30]), .ip2(n1772), .ip3(in2[1]), .ip4(n1064), .op(n833) );
  or2_1 U980 ( .ip1(n2009), .ip2(n833), .op(n836) );
  or2_1 U981 ( .ip1(in1[28]), .ip2(n1058), .op(n832) );
  inv_1 U982 ( .ip(in2[1]), .op(n1058) );
  or2_1 U983 ( .ip1(n1772), .ip2(n1058), .op(n1059) );
  nand2_1 U984 ( .ip1(n832), .ip2(n1059), .op(n834) );
  or2_1 U985 ( .ip1(n834), .ip2(n833), .op(n835) );
  nand2_1 U986 ( .ip1(n836), .ip2(n835), .op(n837) );
  nor2_1 U987 ( .ip1(n837), .ip2(n2024), .op(n850) );
  or2_1 U988 ( .ip1(in1[20]), .ip2(n1058), .op(n838) );
  nand2_1 U989 ( .ip1(n838), .ip2(n1059), .op(n1298) );
  nand2_1 U990 ( .ip1(in1[19]), .ip2(in2[0]), .op(n1296) );
  nand2_1 U991 ( .ip1(n1298), .ip2(n1296), .op(n841) );
  or2_1 U992 ( .ip1(in1[22]), .ip2(in2[1]), .op(n839) );
  nand2_1 U993 ( .ip1(n839), .ip2(n2007), .op(n971) );
  nand2_1 U994 ( .ip1(in2[0]), .ip2(in1[21]), .op(n1937) );
  nand2_1 U995 ( .ip1(n971), .ip2(n1937), .op(n840) );
  nand2_1 U996 ( .ip1(n841), .ip2(n840), .op(n988) );
  nand2_1 U997 ( .ip1(in2[3]), .ip2(n1149), .op(n1815) );
  inv_1 U998 ( .ip(n1815), .op(n2015) );
  nand2_1 U999 ( .ip1(n988), .ip2(n2015), .op(n848) );
  or2_1 U1000 ( .ip1(in1[26]), .ip2(in2[1]), .op(n842) );
  nand2_1 U1001 ( .ip1(n842), .ip2(n2007), .op(n863) );
  nand2_1 U1002 ( .ip1(in1[25]), .ip2(in2[0]), .op(n2006) );
  nand2_1 U1003 ( .ip1(n863), .ip2(n2006), .op(n846) );
  or2_1 U1004 ( .ip1(in1[24]), .ip2(n1058), .op(n843) );
  nand2_1 U1005 ( .ip1(n843), .ip2(n1059), .op(n844) );
  nand2_1 U1006 ( .ip1(in1[23]), .ip2(in2[0]), .op(n1935) );
  nand2_1 U1007 ( .ip1(n844), .ip2(n1935), .op(n845) );
  nand2_1 U1008 ( .ip1(n846), .ip2(n845), .op(n870) );
  nand2_1 U1009 ( .ip1(n2022), .ip2(n870), .op(n847) );
  nand2_1 U1010 ( .ip1(n848), .ip2(n847), .op(n849) );
  not_ab_or_c_or_d U1011 ( .ip1(n987), .ip2(n1946), .ip3(n850), .ip4(n849), 
        .op(n851) );
  nand2_1 U1012 ( .ip1(n2037), .ip2(n851), .op(n852) );
  nand4_1 U1013 ( .ip1(n855), .ip2(n854), .ip3(n853), .ip4(n852), .op(out[30])
         );
  or2_1 U1014 ( .ip1(in2[26]), .ip2(in1[26]), .op(n860) );
  inv_1 U1015 ( .ip(in2[26]), .op(n857) );
  nor2_1 U1016 ( .ip1(in1[26]), .ip2(n857), .op(n1683) );
  inv_1 U1017 ( .ip(in1[26]), .op(n856) );
  nor2_1 U1018 ( .ip1(in2[26]), .ip2(n856), .op(n1601) );
  nor2_1 U1019 ( .ip1(n1683), .ip2(n1601), .op(n1725) );
  nor2_1 U1020 ( .ip1(n1725), .ip2(n1985), .op(n859) );
  nor3_1 U1021 ( .ip1(n1989), .ip2(n857), .ip3(n856), .op(n858) );
  not_ab_or_c_or_d U1022 ( .ip1(n2099), .ip2(n860), .ip3(n859), .ip4(n858), 
        .op(n885) );
  fulladder U1023 ( .a(in1[26]), .b(n862), .ci(n861), .co(n1966), .s(n881) );
  nor2_1 U1024 ( .ip1(n2093), .ip2(n1131), .op(n2075) );
  not_ab_or_c_or_d U1025 ( .ip1(in1[28]), .ip2(n1772), .ip3(n1064), .ip4(n1058), .op(n865) );
  and2_1 U1026 ( .ip1(n863), .ip2(n2009), .op(n864) );
  nor2_1 U1027 ( .ip1(n865), .ip2(n864), .op(n974) );
  nor2_1 U1028 ( .ip1(in2[2]), .ip2(n974), .op(n1479) );
  nand2_1 U1029 ( .ip1(n1509), .ip2(n984), .op(n866) );
  inv_1 U1030 ( .ip(n866), .op(n1478) );
  nor3_1 U1031 ( .ip1(in2[3]), .ip2(n1479), .ip3(n1478), .op(n867) );
  or2_1 U1032 ( .ip1(n2075), .ip2(n867), .op(n1317) );
  inv_1 U1033 ( .ip(n1317), .op(n869) );
  inv_1 U1034 ( .ip(n1198), .op(n2091) );
  nand2_1 U1035 ( .ip1(in2[4]), .ip2(n2093), .op(n868) );
  nand2_1 U1036 ( .ip1(n2091), .ip2(n868), .op(n2077) );
  nor2_1 U1037 ( .ip1(n869), .ip2(n2077), .op(n880) );
  mux2_1 U1038 ( .ip1(n987), .ip2(n989), .s(in2[2]), .op(n1909) );
  nor2_1 U1039 ( .ip1(n1131), .ip2(n1909), .op(n873) );
  inv_1 U1040 ( .ip(n2022), .op(n1941) );
  nor2_1 U1041 ( .ip1(n1941), .ip2(n988), .op(n872) );
  nor2_1 U1042 ( .ip1(n2024), .ip2(n870), .op(n871) );
  nor4_1 U1043 ( .ip1(in2[4]), .ip2(n873), .ip3(n872), .ip4(n871), .op(n878)
         );
  nor2_1 U1044 ( .ip1(n1904), .ip2(n1941), .op(n875) );
  nor2_1 U1045 ( .ip1(n1927), .ip2(n1815), .op(n874) );
  not_ab_or_c_or_d U1046 ( .ip1(n1906), .ip2(n2014), .ip3(n875), .ip4(n874), 
        .op(n1295) );
  inv_1 U1047 ( .ip(n2124), .op(n1978) );
  nor2_1 U1048 ( .ip1(n1295), .ip2(n1978), .op(n876) );
  nor2_1 U1049 ( .ip1(n2037), .ip2(n876), .op(n877) );
  nor2_1 U1050 ( .ip1(n878), .ip2(n877), .op(n879) );
  not_ab_or_c_or_d U1051 ( .ip1(n881), .ip2(n2131), .ip3(n880), .ip4(n879), 
        .op(n884) );
  nor2_1 U1052 ( .ip1(in2[4]), .ip2(in2[3]), .op(n1384) );
  nand2_1 U1053 ( .ip1(n1214), .ip2(n1384), .op(n2027) );
  nor2_1 U1054 ( .ip1(n1875), .ip2(n1149), .op(n882) );
  or2_1 U1055 ( .ip1(n1479), .ip2(n882), .op(n1469) );
  or2_1 U1056 ( .ip1(n2027), .ip2(n1469), .op(n883) );
  nand4_1 U1057 ( .ip1(n885), .ip2(n884), .ip3(n2001), .ip4(n883), .op(out[26]) );
  nand2_1 U1058 ( .ip1(in1[25]), .ip2(n2048), .op(n905) );
  nand2_1 U1059 ( .ip1(in1[26]), .ip2(n2106), .op(n1971) );
  nand2_1 U1060 ( .ip1(n1486), .ip2(in1[28]), .op(n2109) );
  nand2_1 U1061 ( .ip1(in1[27]), .ip2(n1508), .op(n2052) );
  nand4_1 U1062 ( .ip1(n905), .ip2(n1971), .ip3(n2109), .ip4(n2052), .op(n1204) );
  nand2_1 U1063 ( .ip1(n1149), .ip2(n1204), .op(n893) );
  inv_1 U1064 ( .ip(n893), .op(n890) );
  or2_1 U1065 ( .ip1(n886), .ip2(n1149), .op(n888) );
  mux2_1 U1066 ( .ip1(in1[29]), .ip2(in1[30]), .s(in2[0]), .op(n1017) );
  nand2_1 U1067 ( .ip1(n1058), .ip2(n1017), .op(n892) );
  or2_1 U1068 ( .ip1(n892), .ip2(n1149), .op(n887) );
  nand2_1 U1069 ( .ip1(n888), .ip2(n887), .op(n889) );
  nor2_1 U1070 ( .ip1(n890), .ip2(n889), .op(n1522) );
  nand2_1 U1071 ( .ip1(n2091), .ip2(n1384), .op(n1960) );
  nor2_1 U1072 ( .ip1(n1522), .ip2(n1960), .op(n902) );
  nand2_1 U1073 ( .ip1(N316), .ip2(n1508), .op(n891) );
  nand2_1 U1074 ( .ip1(n892), .ip2(n891), .op(n1028) );
  nand2_1 U1075 ( .ip1(n1509), .ip2(n1028), .op(n894) );
  and2_1 U1076 ( .ip1(n894), .ip2(n893), .op(n1521) );
  nor2_1 U1077 ( .ip1(n1521), .ip2(n2027), .op(n901) );
  nor2_1 U1078 ( .ip1(in2[25]), .ip2(in1[25]), .op(n895) );
  nor2_1 U1079 ( .ip1(n895), .ip2(n2046), .op(n900) );
  inv_1 U1080 ( .ip(in1[25]), .op(n896) );
  nor2_1 U1081 ( .ip1(in2[25]), .ip2(n896), .op(n1602) );
  nand2_1 U1082 ( .ip1(in2[25]), .ip2(n896), .op(n1682) );
  inv_1 U1083 ( .ip(n1682), .op(n1541) );
  nor2_1 U1084 ( .ip1(n1602), .ip2(n1541), .op(n1724) );
  or2_1 U1085 ( .ip1(n1724), .ip2(n1985), .op(n898) );
  nand3_1 U1086 ( .ip1(n2092), .ip2(in2[25]), .ip3(in1[25]), .op(n897) );
  nand2_1 U1087 ( .ip1(n898), .ip2(n897), .op(n899) );
  nor4_1 U1088 ( .ip1(n902), .ip2(n901), .ip3(n900), .ip4(n899), .op(n931) );
  inv_1 U1089 ( .ip(n903), .op(n904) );
  nor2_1 U1090 ( .ip1(n1384), .ip2(n904), .op(n955) );
  inv_1 U1091 ( .ip(n955), .op(n1964) );
  nor2_1 U1092 ( .ip1(in2[4]), .ip2(n1815), .op(n2117) );
  nor2_1 U1093 ( .ip1(n1580), .ip2(n2102), .op(n1203) );
  inv_1 U1094 ( .ip(in1[17]), .op(n1306) );
  nor2_1 U1095 ( .ip1(n1306), .ip2(n1782), .op(n1127) );
  nor2_1 U1096 ( .ip1(n1783), .ip2(n1882), .op(n1277) );
  nor2_1 U1097 ( .ip1(n1543), .ip2(n2007), .op(n1191) );
  nor4_1 U1098 ( .ip1(n1203), .ip2(n1127), .ip3(n1277), .ip4(n1191), .op(n1008) );
  nand2_1 U1099 ( .ip1(n2117), .ip2(n1008), .op(n915) );
  nand2_1 U1100 ( .ip1(n1384), .ip2(n1149), .op(n2108) );
  inv_1 U1101 ( .ip(n2108), .op(n2059) );
  inv_1 U1102 ( .ip(in1[23]), .op(n940) );
  nor2_1 U1103 ( .ip1(n940), .ip2(n2102), .op(n1012) );
  inv_1 U1104 ( .ip(n905), .op(n906) );
  inv_1 U1105 ( .ip(in1[22]), .op(n977) );
  nor2_1 U1106 ( .ip1(n1783), .ip2(n977), .op(n1086) );
  inv_1 U1107 ( .ip(in1[24]), .op(n1952) );
  nor2_1 U1108 ( .ip1(n1952), .ip2(n2007), .op(n932) );
  nor4_1 U1109 ( .ip1(n1012), .ip2(n906), .ip3(n1086), .ip4(n932), .op(n2054)
         );
  nand2_1 U1110 ( .ip1(n2059), .ip2(n2054), .op(n914) );
  nor2_1 U1111 ( .ip1(in2[4]), .ip2(n2003), .op(n2119) );
  nand2_1 U1112 ( .ip1(n1508), .ip2(n1359), .op(n910) );
  nand2_1 U1113 ( .ip1(n2048), .ip2(n1554), .op(n909) );
  nand2_1 U1114 ( .ip1(n1486), .ip2(n1391), .op(n908) );
  nand2_1 U1115 ( .ip1(n2106), .ip2(n1661), .op(n907) );
  nand4_1 U1116 ( .ip1(n910), .ip2(n909), .ip3(n908), .ip4(n907), .op(n1133)
         );
  nand2_1 U1117 ( .ip1(n2119), .ip2(n1133), .op(n913) );
  inv_1 U1118 ( .ip(n1384), .op(n911) );
  nor2_1 U1119 ( .ip1(n911), .ip2(n1149), .op(n2115) );
  inv_1 U1120 ( .ip(in1[19]), .op(n1090) );
  nor2_1 U1121 ( .ip1(n1090), .ip2(n2102), .op(n1126) );
  inv_1 U1122 ( .ip(in1[21]), .op(n1002) );
  nor2_1 U1123 ( .ip1(n1002), .ip2(n1782), .op(n1011) );
  inv_1 U1124 ( .ip(in1[18]), .op(n1915) );
  nor2_1 U1125 ( .ip1(n1915), .ip2(n1783), .op(n1190) );
  inv_1 U1126 ( .ip(in1[20]), .op(n1035) );
  nor2_1 U1127 ( .ip1(n1035), .ip2(n2007), .op(n1085) );
  nor4_1 U1128 ( .ip1(n1126), .ip2(n1011), .ip3(n1190), .ip4(n1085), .op(n2060) );
  nand2_1 U1129 ( .ip1(n2115), .ip2(n2060), .op(n912) );
  nand4_1 U1130 ( .ip1(n915), .ip2(n914), .ip3(n913), .ip4(n912), .op(n925) );
  inv_1 U1131 ( .ip(in1[6]), .op(n1407) );
  nand2_1 U1132 ( .ip1(n1486), .ip2(n1407), .op(n1811) );
  nand2_1 U1133 ( .ip1(n1508), .ip2(n1376), .op(n918) );
  nand2_1 U1134 ( .ip1(n2048), .ip2(n1389), .op(n917) );
  inv_1 U1135 ( .ip(in1[8]), .op(n1567) );
  nand2_1 U1136 ( .ip1(n2106), .ip2(n1567), .op(n916) );
  nand4_1 U1137 ( .ip1(n1811), .ip2(n918), .ip3(n917), .ip4(n916), .op(n1007)
         );
  nor2_1 U1138 ( .ip1(n1857), .ip2(n1782), .op(n1505) );
  nor2_1 U1139 ( .ip1(in1[3]), .ip2(in2[0]), .op(n919) );
  not_ab_or_c_or_d U1140 ( .ip1(in2[0]), .ip2(n1472), .ip3(n919), .ip4(n1058), 
        .op(n920) );
  not_ab_or_c_or_d U1141 ( .ip1(n2106), .ip2(in1[4]), .ip3(n1505), .ip4(n920), 
        .op(n1006) );
  mux2_1 U1142 ( .ip1(n1007), .ip2(n1006), .s(in2[2]), .op(n1134) );
  nor2_1 U1143 ( .ip1(in2[3]), .ip2(n1134), .op(n922) );
  nand2_1 U1144 ( .ip1(in2[0]), .ip2(n1770), .op(n1706) );
  inv_1 U1145 ( .ip(in1[1]), .op(n1499) );
  nand2_1 U1146 ( .ip1(n1772), .ip2(n1499), .op(n959) );
  nand3_1 U1147 ( .ip1(n1706), .ip2(n959), .ip3(n1058), .op(n1528) );
  nor2_1 U1148 ( .ip1(n1815), .ip2(n1528), .op(n921) );
  nor2_1 U1149 ( .ip1(n922), .ip2(n921), .op(n1322) );
  nor2_1 U1150 ( .ip1(n1322), .ip2(n1978), .op(n923) );
  nor2_1 U1151 ( .ip1(n2037), .ip2(n923), .op(n924) );
  or2_1 U1152 ( .ip1(n925), .ip2(n924), .op(n930) );
  fulladder U1153 ( .a(in1[25]), .b(n927), .ci(n926), .co(n861), .s(n928) );
  nand2_1 U1154 ( .ip1(n928), .ip2(n2131), .op(n929) );
  nand4_1 U1155 ( .ip1(n931), .ip2(n1964), .ip3(n930), .ip4(n929), .op(out[25]) );
  inv_1 U1156 ( .ip(n932), .op(n933) );
  nand2_1 U1157 ( .ip1(n1486), .ip2(in1[26]), .op(n2050) );
  nand2_1 U1158 ( .ip1(in1[25]), .ip2(n1508), .op(n1970) );
  nand2_1 U1159 ( .ip1(in1[23]), .ip2(n2048), .op(n949) );
  nand4_1 U1160 ( .ip1(n933), .ip2(n2050), .ip3(n1970), .ip4(n949), .op(n1275)
         );
  inv_1 U1161 ( .ip(n1275), .op(n936) );
  nand2_1 U1162 ( .ip1(n1017), .ip2(in2[1]), .op(n934) );
  nand2_1 U1163 ( .ip1(in1[27]), .ip2(n2048), .op(n1969) );
  nand2_1 U1164 ( .ip1(in1[28]), .ip2(n2106), .op(n2049) );
  nand3_1 U1165 ( .ip1(n934), .ip2(n1969), .ip3(n2049), .op(n1256) );
  inv_1 U1166 ( .ip(n1256), .op(n935) );
  mux2_1 U1167 ( .ip1(n936), .ip2(n935), .s(in2[2]), .op(n1400) );
  nor2_1 U1168 ( .ip1(in2[3]), .ip2(n1400), .op(n938) );
  nor2_1 U1169 ( .ip1(n2093), .ip2(n1782), .op(n2105) );
  inv_1 U1170 ( .ip(n2105), .op(n1177) );
  nor2_1 U1171 ( .ip1(n1815), .ip2(n1177), .op(n937) );
  or2_1 U1172 ( .ip1(n938), .ip2(n937), .op(n1381) );
  nor2_1 U1173 ( .ip1(in2[23]), .ip2(in1[23]), .op(n939) );
  nor2_1 U1174 ( .ip1(n939), .ip2(n2046), .op(n944) );
  nor2_1 U1175 ( .ip1(in2[23]), .ip2(n940), .op(n1617) );
  nand2_1 U1176 ( .ip1(in2[23]), .ip2(n940), .op(n1618) );
  inv_1 U1177 ( .ip(n1618), .op(n1612) );
  nor2_1 U1178 ( .ip1(n1617), .ip2(n1612), .op(n1719) );
  or2_1 U1179 ( .ip1(n1719), .ip2(n1985), .op(n942) );
  nand3_1 U1180 ( .ip1(n2092), .ip2(in2[23]), .ip3(in1[23]), .op(n941) );
  nand2_1 U1181 ( .ip1(n942), .ip2(n941), .op(n943) );
  not_ab_or_c_or_d U1182 ( .ip1(n2098), .ip2(n1381), .ip3(n944), .ip4(n943), 
        .op(n968) );
  nand2_1 U1183 ( .ip1(n1508), .ip2(n1389), .op(n948) );
  nand2_1 U1184 ( .ip1(n2048), .ip2(n1359), .op(n947) );
  nand2_1 U1185 ( .ip1(n1486), .ip2(n1567), .op(n946) );
  nand2_1 U1186 ( .ip1(n2106), .ip2(n1391), .op(n945) );
  nand4_1 U1187 ( .ip1(n948), .ip2(n947), .ip3(n946), .ip4(n945), .op(n1259)
         );
  inv_1 U1188 ( .ip(n1259), .op(n1099) );
  nand2_1 U1189 ( .ip1(n1946), .ip2(n1099), .op(n953) );
  nand2_1 U1190 ( .ip1(in1[17]), .ip2(n1508), .op(n1188) );
  nand2_1 U1191 ( .ip1(in1[19]), .ip2(n2048), .op(n1082) );
  nand2_1 U1192 ( .ip1(n1486), .ip2(in1[16]), .op(n1200) );
  nand2_1 U1193 ( .ip1(in1[18]), .ip2(n2106), .op(n1129) );
  nand4_1 U1194 ( .ip1(n1188), .ip2(n1082), .ip3(n1200), .ip4(n1129), .op(
        n2118) );
  nand2_1 U1195 ( .ip1(n2022), .ip2(n2118), .op(n952) );
  nand2_1 U1196 ( .ip1(in1[13]), .ip2(n1508), .op(n1278) );
  nand2_1 U1197 ( .ip1(in1[15]), .ip2(n2048), .op(n1187) );
  nand2_1 U1198 ( .ip1(n1486), .ip2(in1[12]), .op(n1337) );
  nand2_1 U1199 ( .ip1(in1[14]), .ip2(n2106), .op(n1201) );
  nand4_1 U1200 ( .ip1(n1278), .ip2(n1187), .ip3(n1337), .ip4(n1201), .op(
        n1972) );
  nand2_1 U1201 ( .ip1(n2015), .ip2(n1972), .op(n951) );
  nand2_1 U1202 ( .ip1(in1[21]), .ip2(n1508), .op(n1083) );
  nand2_1 U1203 ( .ip1(n1486), .ip2(in1[20]), .op(n1128) );
  nand2_1 U1204 ( .ip1(in1[22]), .ip2(n2106), .op(n1013) );
  nand4_1 U1205 ( .ip1(n1083), .ip2(n949), .ip3(n1128), .ip4(n1013), .op(n2116) );
  nand2_1 U1206 ( .ip1(n2014), .ip2(n2116), .op(n950) );
  nand4_1 U1207 ( .ip1(n953), .ip2(n952), .ip3(n951), .ip4(n950), .op(n956) );
  nor2_1 U1208 ( .ip1(n1400), .ip2(n1960), .op(n954) );
  not_ab_or_c_or_d U1209 ( .ip1(n2037), .ip2(n956), .ip3(n955), .ip4(n954), 
        .op(n967) );
  nand2_1 U1210 ( .ip1(n1508), .ip2(n1857), .op(n1810) );
  nand2_1 U1211 ( .ip1(n2048), .ip2(n1376), .op(n958) );
  inv_1 U1212 ( .ip(in1[4]), .op(n1807) );
  nand2_1 U1213 ( .ip1(n1486), .ip2(n1807), .op(n1510) );
  nand2_1 U1214 ( .ip1(n2106), .ip2(n1407), .op(n957) );
  nand4_1 U1215 ( .ip1(n1810), .ip2(n958), .ip3(n1510), .ip4(n957), .op(n1260)
         );
  nor2_1 U1216 ( .ip1(n1472), .ip2(n2007), .op(n961) );
  and3_1 U1217 ( .ip1(in2[1]), .ip2(n1706), .ip3(n959), .op(n960) );
  not_ab_or_c_or_d U1218 ( .ip1(n2048), .ip2(in1[3]), .ip3(n961), .ip4(n960), 
        .op(n1806) );
  mux2_1 U1219 ( .ip1(n1260), .ip2(n1806), .s(in2[2]), .op(n1385) );
  inv_1 U1220 ( .ip(in2[3]), .op(n1131) );
  nand2_1 U1221 ( .ip1(in2[4]), .ip2(n1131), .op(n1199) );
  inv_1 U1222 ( .ip(n1199), .op(n1213) );
  nand2_1 U1223 ( .ip1(n2124), .ip2(n1213), .op(n1150) );
  or2_1 U1224 ( .ip1(n1385), .ip2(n1150), .op(n966) );
  fulladder U1225 ( .a(in1[23]), .b(n963), .ci(n962), .co(n1933), .s(n964) );
  nand2_1 U1226 ( .ip1(n964), .ip2(n2131), .op(n965) );
  nand4_1 U1227 ( .ip1(n968), .ip2(n967), .ip3(n966), .ip4(n965), .op(out[23])
         );
  or2_1 U1228 ( .ip1(in2[22]), .ip2(in1[22]), .op(n982) );
  nor2_1 U1229 ( .ip1(n1406), .ip2(n1150), .op(n981) );
  nand2_1 U1230 ( .ip1(n2015), .ip2(n1875), .op(n975) );
  inv_1 U1231 ( .ip(n2006), .op(n969) );
  not_ab_or_c_or_d U1232 ( .ip1(in1[24]), .ip2(n1772), .ip3(n969), .ip4(n1058), 
        .op(n970) );
  or2_1 U1233 ( .ip1(n1935), .ip2(n970), .op(n973) );
  or2_1 U1234 ( .ip1(n971), .ip2(n970), .op(n972) );
  nand2_1 U1235 ( .ip1(n973), .ip2(n972), .op(n1468) );
  mux2_1 U1236 ( .ip1(n1468), .ip2(n974), .s(n1509), .op(n1887) );
  nand2_1 U1237 ( .ip1(n1131), .ip2(n1887), .op(n983) );
  nand2_1 U1238 ( .ip1(n975), .ip2(n983), .op(n1409) );
  inv_1 U1239 ( .ip(in2[22]), .op(n976) );
  nor2_1 U1240 ( .ip1(n976), .ip2(in1[22]), .op(n1611) );
  nor2_1 U1241 ( .ip1(in2[22]), .ip2(n977), .op(n1619) );
  nor2_1 U1242 ( .ip1(n1611), .ip2(n1619), .op(n1718) );
  nor2_1 U1243 ( .ip1(n1718), .ip2(n1985), .op(n979) );
  nor3_1 U1244 ( .ip1(n1989), .ip2(n977), .ip3(n976), .op(n978) );
  ab_or_c_or_d U1245 ( .ip1(n2098), .ip2(n1409), .ip3(n979), .ip4(n978), .op(
        n980) );
  not_ab_or_c_or_d U1246 ( .ip1(n2099), .ip2(n982), .ip3(n981), .ip4(n980), 
        .op(n1000) );
  inv_1 U1247 ( .ip(n983), .op(n986) );
  nor2_1 U1248 ( .ip1(N316), .ip2(n1149), .op(n1257) );
  not_ab_or_c_or_d U1249 ( .ip1(n984), .ip2(n1149), .ip3(n1257), .ip4(n1131), 
        .op(n985) );
  nor2_1 U1250 ( .ip1(n986), .ip2(n985), .op(n1428) );
  nor2_1 U1251 ( .ip1(n1428), .ip2(n2077), .op(n994) );
  mux2_1 U1252 ( .ip1(n988), .ip2(n987), .s(in2[2]), .op(n992) );
  nor2_1 U1253 ( .ip1(n989), .ip2(n1509), .op(n990) );
  not_ab_or_c_or_d U1254 ( .ip1(in2[2]), .ip2(n1906), .ip3(n1131), .ip4(n990), 
        .op(n991) );
  not_ab_or_c_or_d U1255 ( .ip1(n992), .ip2(n1131), .ip3(n991), .ip4(n1907), 
        .op(n993) );
  nor2_1 U1256 ( .ip1(n994), .ip2(n993), .op(n999) );
  fulladder U1257 ( .a(in1[22]), .b(n996), .ci(n995), .co(n962), .s(n997) );
  nand2_1 U1258 ( .ip1(n997), .ip2(n2131), .op(n998) );
  nand4_1 U1259 ( .ip1(n1000), .ip2(n999), .ip3(n2001), .ip4(n998), .op(
        out[22]) );
  or2_1 U1260 ( .ip1(in2[21]), .ip2(in1[21]), .op(n1005) );
  inv_1 U1261 ( .ip(in2[21]), .op(n1001) );
  nor2_1 U1262 ( .ip1(in1[21]), .ip2(n1001), .op(n1613) );
  nor2_1 U1263 ( .ip1(in2[21]), .ip2(n1002), .op(n1553) );
  nor2_1 U1264 ( .ip1(n1613), .ip2(n1553), .op(n1717) );
  nor2_1 U1265 ( .ip1(n1717), .ip2(n1985), .op(n1004) );
  nor3_1 U1266 ( .ip1(n1989), .ip2(n1002), .ip3(n1001), .op(n1003) );
  not_ab_or_c_or_d U1267 ( .ip1(n2099), .ip2(n1005), .ip3(n1004), .ip4(n1003), 
        .op(n1033) );
  inv_1 U1268 ( .ip(n1150), .op(n1103) );
  mux2_1 U1269 ( .ip1(n1006), .ip2(n1528), .s(in2[2]), .op(n1841) );
  inv_1 U1270 ( .ip(n1841), .op(n1024) );
  mux2_1 U1271 ( .ip1(n1133), .ip2(n1007), .s(in2[2]), .op(n1222) );
  inv_1 U1272 ( .ip(n1008), .op(n2062) );
  nor2_1 U1273 ( .ip1(n2060), .ip2(n1509), .op(n1009) );
  not_ab_or_c_or_d U1274 ( .ip1(in2[2]), .ip2(n2062), .ip3(in2[3]), .ip4(n1009), .op(n1010) );
  not_ab_or_c_or_d U1275 ( .ip1(n1222), .ip2(in2[3]), .ip3(n1010), .ip4(n1907), 
        .op(n1023) );
  nor2_1 U1276 ( .ip1(n1012), .ip2(n1011), .op(n1014) );
  nand2_1 U1277 ( .ip1(in1[24]), .ip2(n1486), .op(n1968) );
  nand3_1 U1278 ( .ip1(n1014), .ip2(n1968), .ip3(n1013), .op(n1205) );
  mux2_1 U1279 ( .ip1(n1205), .ip2(n1204), .s(in2[2]), .op(n1015) );
  nor2_1 U1280 ( .ip1(in2[3]), .ip2(n1015), .op(n1847) );
  or2_1 U1281 ( .ip1(in2[3]), .ip2(n1847), .op(n1019) );
  nand2_1 U1282 ( .ip1(n1149), .ip2(n1058), .op(n1016) );
  mux2_1 U1283 ( .ip1(n1017), .ip2(N316), .s(n1016), .op(n2076) );
  inv_1 U1284 ( .ip(n2076), .op(n1842) );
  or2_1 U1285 ( .ip1(n1842), .ip2(n1847), .op(n1018) );
  nand2_1 U1286 ( .ip1(n1019), .ip2(n1018), .op(n1020) );
  nor2_1 U1287 ( .ip1(in2[4]), .ip2(n1020), .op(n1021) );
  nor2_1 U1288 ( .ip1(n1021), .ip2(n2077), .op(n1022) );
  not_ab_or_c_or_d U1289 ( .ip1(n1103), .ip2(n1024), .ip3(n1023), .ip4(n1022), 
        .op(n1032) );
  fulladder U1290 ( .a(in1[21]), .b(n1026), .ci(n1025), .co(n995), .s(n1027)
         );
  nand2_1 U1291 ( .ip1(n1027), .ip2(n2131), .op(n1031) );
  inv_1 U1292 ( .ip(in2[2]), .op(n1149) );
  nand2_1 U1293 ( .ip1(n1028), .ip2(n1149), .op(n1215) );
  inv_1 U1294 ( .ip(n1215), .op(n2073) );
  nor2_1 U1295 ( .ip1(n2073), .ip2(n1131), .op(n1029) );
  nor2_1 U1296 ( .ip1(n1847), .ip2(n1029), .op(n1865) );
  nand2_1 U1297 ( .ip1(n2098), .ip2(n1865), .op(n1030) );
  nand4_1 U1298 ( .ip1(n1033), .ip2(n1032), .ip3(n1031), .ip4(n1030), .op(
        out[21]) );
  or2_1 U1299 ( .ip1(in2[20]), .ip2(in1[20]), .op(n1038) );
  inv_1 U1300 ( .ip(in2[20]), .op(n1034) );
  nor2_1 U1301 ( .ip1(in1[20]), .ip2(n1034), .op(n1610) );
  nor2_1 U1302 ( .ip1(in2[20]), .ip2(n1035), .op(n1552) );
  nor2_1 U1303 ( .ip1(n1610), .ip2(n1552), .op(n1716) );
  nor2_1 U1304 ( .ip1(n1716), .ip2(n1985), .op(n1037) );
  nor3_1 U1305 ( .ip1(n1989), .ip2(n1035), .ip3(n1034), .op(n1036) );
  not_ab_or_c_or_d U1306 ( .ip1(n2099), .ip2(n1038), .ip3(n1037), .ip4(n1036), 
        .op(n1080) );
  fulladder U1307 ( .a(in1[20]), .b(n1040), .ci(n1039), .co(n1025), .s(n1074)
         );
  nor2_1 U1308 ( .ip1(n1407), .ip2(n2102), .op(n1439) );
  nor2_1 U1309 ( .ip1(n1567), .ip2(n1782), .op(n1362) );
  not_ab_or_c_or_d U1310 ( .ip1(n1486), .ip2(in1[5]), .ip3(n1439), .ip4(n1362), 
        .op(n1041) );
  nand2_1 U1311 ( .ip1(in1[7]), .ip2(n2106), .op(n1419) );
  nand2_1 U1312 ( .ip1(n1041), .ip2(n1419), .op(n1350) );
  nor2_1 U1313 ( .ip1(n2003), .ip2(n1350), .op(n1053) );
  nor2_1 U1314 ( .ip1(in1[14]), .ip2(n2102), .op(n1043) );
  nor2_1 U1315 ( .ip1(in1[13]), .ip2(n1783), .op(n1042) );
  not_ab_or_c_or_d U1316 ( .ip1(n1044), .ip2(n1058), .ip3(n1043), .ip4(n1042), 
        .op(n2004) );
  or2_1 U1317 ( .ip1(in1[18]), .ip2(n1058), .op(n1045) );
  nand2_1 U1318 ( .ip1(n1045), .ip2(n1059), .op(n1151) );
  nand2_1 U1319 ( .ip1(n1151), .ip2(n1153), .op(n1048) );
  or2_1 U1320 ( .ip1(in1[20]), .ip2(in2[1]), .op(n1046) );
  nand2_1 U1321 ( .ip1(n1046), .ip2(n2007), .op(n1055) );
  nand2_1 U1322 ( .ip1(n1296), .ip2(n1055), .op(n1047) );
  nand2_1 U1323 ( .ip1(n1048), .ip2(n1047), .op(n2016) );
  nor2_1 U1324 ( .ip1(n2016), .ip2(n1509), .op(n1049) );
  not_ab_or_c_or_d U1325 ( .ip1(in2[2]), .ip2(n2004), .ip3(in2[3]), .ip4(n1049), .op(n1052) );
  nor2_1 U1326 ( .ip1(n1661), .ip2(n1782), .op(n1232) );
  nor2_1 U1327 ( .ip1(n1391), .ip2(n2102), .op(n1361) );
  nand2_1 U1328 ( .ip1(n1486), .ip2(in1[9]), .op(n1416) );
  inv_1 U1329 ( .ip(n1416), .op(n1050) );
  nor2_1 U1330 ( .ip1(n1359), .ip2(n2007), .op(n1303) );
  nor4_1 U1331 ( .ip1(n1232), .ip2(n1361), .ip3(n1050), .ip4(n1303), .op(n1237) );
  inv_1 U1332 ( .ip(n1237), .op(n1945) );
  nor2_1 U1333 ( .ip1(n1815), .ip2(n1945), .op(n1051) );
  nor4_1 U1334 ( .ip1(n1053), .ip2(n1052), .ip3(n1051), .ip4(n1907), .op(n1073) );
  or2_1 U1335 ( .ip1(in1[22]), .ip2(n1058), .op(n1054) );
  nand2_1 U1336 ( .ip1(n1054), .ip2(n1059), .op(n1938) );
  nand2_1 U1337 ( .ip1(n1938), .ip2(n1935), .op(n1057) );
  nand2_1 U1338 ( .ip1(n1055), .ip2(n1937), .op(n1056) );
  nand2_1 U1339 ( .ip1(n1057), .ip2(n1056), .op(n1156) );
  or2_1 U1340 ( .ip1(in1[26]), .ip2(n1058), .op(n1060) );
  nand2_1 U1341 ( .ip1(n1060), .ip2(n1059), .op(n2005) );
  nand2_1 U1342 ( .ip1(n2005), .ip2(n2009), .op(n1063) );
  or2_1 U1343 ( .ip1(in1[24]), .ip2(in2[1]), .op(n1061) );
  nand2_1 U1344 ( .ip1(n1061), .ip2(n2007), .op(n1936) );
  nand2_1 U1345 ( .ip1(n1936), .ip2(n2006), .op(n1062) );
  nand2_1 U1346 ( .ip1(n1063), .ip2(n1062), .op(n1157) );
  mux2_1 U1347 ( .ip1(n1156), .ip2(n1157), .s(in2[2]), .op(n1233) );
  and2_1 U1348 ( .ip1(n1131), .ip2(n1233), .op(n1452) );
  nor2_1 U1349 ( .ip1(n2093), .ip2(n1149), .op(n1107) );
  nor2_1 U1350 ( .ip1(in1[30]), .ip2(n2102), .op(n1066) );
  not_ab_or_c_or_d U1351 ( .ip1(in1[28]), .ip2(n1772), .ip3(in2[1]), .ip4(
        n1064), .op(n1065) );
  ab_or_c_or_d U1352 ( .ip1(n1486), .ip2(n2093), .ip3(n1066), .ip4(n1065), 
        .op(n1229) );
  nor2_1 U1353 ( .ip1(n1509), .ip2(n1229), .op(n2028) );
  or2_1 U1354 ( .ip1(n2028), .ip2(n1131), .op(n1068) );
  nor2_1 U1355 ( .ip1(n1107), .ip2(n1068), .op(n1447) );
  inv_1 U1356 ( .ip(n1922), .op(n1067) );
  nor2_1 U1357 ( .ip1(n1447), .ip2(n1067), .op(n1070) );
  inv_1 U1358 ( .ip(n1068), .op(n1448) );
  inv_1 U1359 ( .ip(n2098), .op(n1912) );
  nor2_1 U1360 ( .ip1(n1448), .ip2(n1912), .op(n1069) );
  nor2_1 U1361 ( .ip1(n1070), .ip2(n1069), .op(n1071) );
  nor2_1 U1362 ( .ip1(n1452), .ip2(n1071), .op(n1072) );
  not_ab_or_c_or_d U1363 ( .ip1(n1074), .ip2(n2131), .ip3(n1073), .ip4(n1072), 
        .op(n1079) );
  nor2_1 U1364 ( .ip1(n1807), .ip2(n1782), .op(n1440) );
  nor2_1 U1365 ( .ip1(in1[2]), .ip2(in2[0]), .op(n1075) );
  not_ab_or_c_or_d U1366 ( .ip1(in2[0]), .ip2(n1499), .ip3(n1075), .ip4(n1058), 
        .op(n1076) );
  not_ab_or_c_or_d U1367 ( .ip1(n2106), .ip2(in1[3]), .ip3(n1440), .ip4(n1076), 
        .op(n1347) );
  nand2_1 U1368 ( .ip1(in1[0]), .ip2(n2048), .op(n1077) );
  mux2_1 U1369 ( .ip1(n1347), .ip2(n1077), .s(n1509), .op(n1458) );
  or2_1 U1370 ( .ip1(n1458), .ip2(n1150), .op(n1078) );
  nand4_1 U1371 ( .ip1(n1080), .ip2(n1079), .ip3(n2001), .ip4(n1078), .op(
        out[20]) );
  nor2_1 U1372 ( .ip1(in1[19]), .ip2(in2[19]), .op(n1081) );
  nor2_1 U1373 ( .ip1(n1081), .ip2(n2046), .op(n1095) );
  nand2_1 U1374 ( .ip1(in2[19]), .ip2(n1090), .op(n1608) );
  inv_1 U1375 ( .ip(n1608), .op(n1620) );
  nor2_1 U1376 ( .ip1(in2[19]), .ip2(n1090), .op(n1606) );
  nor2_1 U1377 ( .ip1(n1620), .ip2(n1606), .op(n1734) );
  nor2_1 U1378 ( .ip1(n1734), .ip2(n1985), .op(n1094) );
  nand2_1 U1379 ( .ip1(n1083), .ip2(n1082), .op(n1084) );
  nor3_1 U1380 ( .ip1(n1086), .ip2(n1085), .ip3(n1084), .op(n1394) );
  nor2_1 U1381 ( .ip1(n1394), .ip2(n1509), .op(n1087) );
  not_ab_or_c_or_d U1382 ( .ip1(in2[2]), .ip2(n1275), .ip3(in2[3]), .ip4(n1087), .op(n1109) );
  inv_1 U1383 ( .ip(n1109), .op(n1089) );
  mux2_1 U1384 ( .ip1(n1256), .ip2(n2105), .s(in2[2]), .op(n1265) );
  or2_1 U1385 ( .ip1(n1265), .ip2(n1131), .op(n1088) );
  nand2_1 U1386 ( .ip1(n1089), .ip2(n1088), .op(n1822) );
  nor2_1 U1387 ( .ip1(n1822), .ip2(n1912), .op(n1093) );
  inv_1 U1388 ( .ip(in2[19]), .op(n1091) );
  nor3_1 U1389 ( .ip1(n1989), .ip2(n1091), .ip3(n1090), .op(n1092) );
  nor4_1 U1390 ( .ip1(n1095), .ip2(n1094), .ip3(n1093), .ip4(n1092), .op(n1112) );
  fulladder U1391 ( .a(in1[19]), .b(n1097), .ci(n1096), .co(n1039), .s(n1106)
         );
  nor2_1 U1392 ( .ip1(n1260), .ip2(n1149), .op(n1098) );
  not_ab_or_c_or_d U1393 ( .ip1(n1099), .ip2(n1149), .ip3(n1131), .ip4(n1098), 
        .op(n1102) );
  nor2_1 U1394 ( .ip1(n2118), .ip2(n2024), .op(n1101) );
  nor2_1 U1395 ( .ip1(n1941), .ip2(n1972), .op(n1100) );
  nor4_1 U1396 ( .ip1(n1102), .ip2(n1101), .ip3(n1100), .ip4(n1907), .op(n1105) );
  nand2_1 U1397 ( .ip1(n1103), .ip2(n1149), .op(n1926) );
  nor2_1 U1398 ( .ip1(n1806), .ip2(n1926), .op(n1104) );
  not_ab_or_c_or_d U1399 ( .ip1(n1106), .ip2(n2131), .ip3(n1105), .ip4(n1104), 
        .op(n1111) );
  not_ab_or_c_or_d U1400 ( .ip1(n1149), .ip2(n1256), .ip3(n1107), .ip4(n1131), 
        .op(n1108) );
  nor2_1 U1401 ( .ip1(n1109), .ip2(n1108), .op(n1829) );
  nand2_1 U1402 ( .ip1(n1922), .ip2(n1829), .op(n1110) );
  nand4_1 U1403 ( .ip1(n1112), .ip2(n1111), .ip3(n2001), .ip4(n1110), .op(
        out[19]) );
  nand2_1 U1404 ( .ip1(in2[17]), .ip2(n1306), .op(n1674) );
  inv_1 U1405 ( .ip(in2[17]), .op(n1113) );
  nand2_1 U1406 ( .ip1(in1[17]), .ip2(n1113), .op(n1605) );
  and2_1 U1407 ( .ip1(n1674), .ip2(n1605), .op(n1733) );
  nor2_1 U1408 ( .ip1(n1733), .ip2(n1985), .op(n1121) );
  nor3_1 U1409 ( .ip1(n1989), .ip2(n1306), .ip3(n1113), .op(n1120) );
  nor2_1 U1410 ( .ip1(n1522), .ip2(n2077), .op(n1115) );
  nor2_1 U1411 ( .ip1(n1521), .ip2(n1912), .op(n1114) );
  nor2_1 U1412 ( .ip1(n1115), .ip2(n1114), .op(n1116) );
  nor2_1 U1413 ( .ip1(n1116), .ip2(n1131), .op(n1119) );
  nor2_1 U1414 ( .ip1(in1[17]), .ip2(in2[17]), .op(n1117) );
  nor2_1 U1415 ( .ip1(n1117), .ip2(n2046), .op(n1118) );
  nor4_1 U1416 ( .ip1(n1121), .ip2(n1120), .ip3(n1119), .ip4(n1118), .op(n1141) );
  fulladder U1417 ( .a(in1[17]), .b(n1123), .ci(n1122), .co(n1924), .s(n1125)
         );
  nor2_1 U1418 ( .ip1(n1528), .ip2(n1926), .op(n1124) );
  inv_1 U1419 ( .ip(n2001), .op(n1928) );
  not_ab_or_c_or_d U1420 ( .ip1(n1125), .ip2(n2131), .ip3(n1124), .ip4(n1928), 
        .op(n1140) );
  inv_1 U1421 ( .ip(n2077), .op(n1999) );
  nor2_1 U1422 ( .ip1(n2098), .ip2(n1999), .op(n1132) );
  nor2_1 U1423 ( .ip1(n1127), .ip2(n1126), .op(n1130) );
  nand3_1 U1424 ( .ip1(n1130), .ip2(n1129), .ip3(n1128), .op(n1849) );
  mux2_1 U1425 ( .ip1(n1849), .ip2(n1205), .s(n1509), .op(n1333) );
  nand2_1 U1426 ( .ip1(n1333), .ip2(n1131), .op(n1516) );
  or2_1 U1427 ( .ip1(n1132), .ip2(n1516), .op(n1139) );
  nand2_1 U1428 ( .ip1(n2022), .ip2(n1133), .op(n1137) );
  or2_1 U1429 ( .ip1(n2062), .ip2(n2024), .op(n1136) );
  nand2_1 U1430 ( .ip1(in2[3]), .ip2(n1134), .op(n1135) );
  nand4_1 U1431 ( .ip1(n2037), .ip2(n1137), .ip3(n1136), .ip4(n1135), .op(
        n1138) );
  nand4_1 U1432 ( .ip1(n1141), .ip2(n1140), .ip3(n1139), .ip4(n1138), .op(
        out[17]) );
  or2_1 U1433 ( .ip1(in2[16]), .ip2(in1[16]), .op(n1146) );
  nand2_1 U1434 ( .ip1(in2[16]), .ip2(n1543), .op(n1675) );
  inv_1 U1435 ( .ip(n1675), .op(n1142) );
  nor2_1 U1436 ( .ip1(in2[16]), .ip2(n1543), .op(n1603) );
  nor2_1 U1437 ( .ip1(n1142), .ip2(n1603), .op(n1732) );
  nor2_1 U1438 ( .ip1(n1732), .ip2(n1985), .op(n1145) );
  inv_1 U1439 ( .ip(in2[16]), .op(n1143) );
  nor3_1 U1440 ( .ip1(n1989), .ip2(n1143), .ip3(n1543), .op(n1144) );
  not_ab_or_c_or_d U1441 ( .ip1(n2099), .ip2(n1146), .ip3(n1145), .ip4(n1144), 
        .op(n1170) );
  fulladder U1442 ( .a(in1[16]), .b(n1148), .ci(n1147), .co(n1122), .s(n1163)
         );
  nand3_1 U1443 ( .ip1(in1[0]), .ip2(n2048), .ip3(n1149), .op(n1769) );
  nor2_1 U1444 ( .ip1(n1769), .ip2(n1150), .op(n1162) );
  nand2_1 U1445 ( .ip1(n1296), .ip2(n1151), .op(n1155) );
  nand2_1 U1446 ( .ip1(in1[16]), .ip2(n1772), .op(n1152) );
  nand3_1 U1447 ( .ip1(n1153), .ip2(n1152), .ip3(n1058), .op(n1154) );
  nand2_1 U1448 ( .ip1(n1155), .ip2(n1154), .op(n1438) );
  mux2_1 U1449 ( .ip1(n1438), .ip2(n1156), .s(in2[2]), .op(n1793) );
  inv_1 U1450 ( .ip(n1157), .op(n1159) );
  inv_1 U1451 ( .ip(n1229), .op(n1158) );
  mux2_1 U1452 ( .ip1(n1159), .ip2(n1158), .s(in2[2]), .op(n1962) );
  nor2_1 U1453 ( .ip1(n1962), .ip2(n1131), .op(n1160) );
  or2_1 U1454 ( .ip1(n2091), .ip2(n1214), .op(n1798) );
  nand2_1 U1455 ( .ip1(n2100), .ip2(n1798), .op(n1854) );
  not_ab_or_c_or_d U1456 ( .ip1(n1793), .ip2(n1131), .ip3(n1160), .ip4(n1854), 
        .op(n1161) );
  not_ab_or_c_or_d U1457 ( .ip1(n1163), .ip2(n2131), .ip3(n1162), .ip4(n1161), 
        .op(n1169) );
  nor2_1 U1458 ( .ip1(n2004), .ip2(n1509), .op(n1164) );
  not_ab_or_c_or_d U1459 ( .ip1(in2[2]), .ip2(n1237), .ip3(in2[3]), .ip4(n1164), .op(n1166) );
  nor2_1 U1460 ( .ip1(n1347), .ip2(n2003), .op(n1165) );
  not_ab_or_c_or_d U1461 ( .ip1(n1350), .ip2(n2015), .ip3(n1166), .ip4(n1165), 
        .op(n1167) );
  or2_1 U1462 ( .ip1(n1167), .ip2(n1907), .op(n1168) );
  nand4_1 U1463 ( .ip1(n1170), .ip2(n1169), .ip3(n2001), .ip4(n1168), .op(
        out[16]) );
  nor2_1 U1464 ( .ip1(n1131), .ip2(n1385), .op(n1172) );
  nor2_1 U1465 ( .ip1(n1941), .ip2(n1259), .op(n1171) );
  not_ab_or_c_or_d U1466 ( .ip1(n1972), .ip2(n2014), .ip3(n1172), .ip4(n1171), 
        .op(n2101) );
  nor2_1 U1467 ( .ip1(n2101), .ip2(n1907), .op(n1183) );
  nor2_1 U1468 ( .ip1(in2[15]), .ip2(n1580), .op(n1574) );
  inv_1 U1469 ( .ip(n1574), .op(n1672) );
  nor2_1 U1470 ( .ip1(n1985), .ip2(n1672), .op(n1182) );
  nor2_1 U1471 ( .ip1(in1[15]), .ip2(n1748), .op(n1175) );
  nor2_1 U1472 ( .ip1(op[1]), .ip2(n1580), .op(n1174) );
  inv_1 U1473 ( .ip(in2[15]), .op(n1173) );
  nor4_1 U1474 ( .ip1(n1176), .ip2(n1175), .ip3(n1174), .ip4(n1173), .op(n1181) );
  nand2_1 U1475 ( .ip1(n2099), .ip2(in1[15]), .op(n1179) );
  nand2_1 U1476 ( .ip1(in2[4]), .ip2(n1214), .op(n1821) );
  inv_1 U1477 ( .ip(n1821), .op(n1876) );
  nor2_1 U1478 ( .ip1(n2024), .ip2(n1177), .op(n2097) );
  nand2_1 U1479 ( .ip1(n1876), .ip2(n2097), .op(n1178) );
  nand2_1 U1480 ( .ip1(n1179), .ip2(n1178), .op(n1180) );
  nor4_1 U1481 ( .ip1(n1183), .ip2(n1182), .ip3(n1181), .ip4(n1180), .op(n1197) );
  fulladder U1482 ( .a(in1[15]), .b(n1185), .ci(n1184), .co(n1147), .s(n1186)
         );
  nand2_1 U1483 ( .ip1(n1186), .ip2(n2131), .op(n1196) );
  inv_1 U1484 ( .ip(n1854), .op(n1893) );
  nand2_1 U1485 ( .ip1(n1188), .ip2(n1187), .op(n1189) );
  nor3_1 U1486 ( .ip1(n1191), .ip2(n1190), .ip3(n1189), .op(n1813) );
  nand2_1 U1487 ( .ip1(n2014), .ip2(n1813), .op(n1194) );
  nand2_1 U1488 ( .ip1(in2[3]), .ip2(n1400), .op(n1193) );
  nand2_1 U1489 ( .ip1(n2022), .ip2(n1394), .op(n1192) );
  nand4_1 U1490 ( .ip1(n1893), .ip2(n1194), .ip3(n1193), .ip4(n1192), .op(
        n1195) );
  nand4_1 U1491 ( .ip1(n1197), .ip2(n2001), .ip3(n1196), .ip4(n1195), .op(
        out[15]) );
  nor2_1 U1492 ( .ip1(n1199), .ip2(n1198), .op(n1845) );
  nand2_1 U1493 ( .ip1(n1201), .ip2(n1200), .op(n1202) );
  not_ab_or_c_or_d U1494 ( .ip1(n2048), .ip2(in1[13]), .ip3(n1203), .ip4(n1202), .op(n1852) );
  inv_1 U1495 ( .ip(n1204), .op(n1208) );
  nor2_1 U1496 ( .ip1(n1941), .ip2(n1849), .op(n1207) );
  nor2_1 U1497 ( .ip1(n1815), .ip2(n1205), .op(n1206) );
  ab_or_c_or_d U1498 ( .ip1(n1946), .ip2(n1208), .ip3(n1207), .ip4(n1206), 
        .op(n1209) );
  not_ab_or_c_or_d U1499 ( .ip1(n1852), .ip2(n2014), .ip3(n1854), .ip4(n1209), 
        .op(n1221) );
  nor2_1 U1500 ( .ip1(n2046), .ip2(n1554), .op(n1219) );
  inv_1 U1501 ( .ip(in2[13]), .op(n1211) );
  nand2_1 U1502 ( .ip1(in1[13]), .ip2(n1211), .op(n1623) );
  nor2_1 U1503 ( .ip1(n1623), .ip2(n1985), .op(n1218) );
  nor2_1 U1504 ( .ip1(n1985), .ip2(in1[13]), .op(n1210) );
  not_ab_or_c_or_d U1505 ( .ip1(in1[13]), .ip2(n2092), .ip3(n2099), .ip4(n1210), .op(n1212) );
  nor2_1 U1506 ( .ip1(n1212), .ip2(n1211), .op(n1217) );
  nand2_1 U1507 ( .ip1(n1214), .ip2(n1213), .op(n1324) );
  nor2_1 U1508 ( .ip1(n1215), .ip2(n1324), .op(n1216) );
  or4_1 U1509 ( .ip1(n1219), .ip2(n1218), .ip3(n1217), .ip4(n1216), .op(n1220)
         );
  not_ab_or_c_or_d U1510 ( .ip1(n2076), .ip2(n1845), .ip3(n1221), .ip4(n1220), 
        .op(n1228) );
  mux2_1 U1511 ( .ip1(n1222), .ip2(n1841), .s(in2[3]), .op(n2055) );
  or2_1 U1512 ( .ip1(n2055), .ip2(n1907), .op(n1227) );
  nand2_1 U1513 ( .ip1(n1874), .ip2(n2075), .op(n1373) );
  fulladder U1514 ( .a(in1[13]), .b(n1224), .ci(n1223), .co(n1894), .s(n1225)
         );
  nand2_1 U1515 ( .ip1(n1225), .ip2(n2131), .op(n1226) );
  nand4_1 U1516 ( .ip1(n1228), .ip2(n1227), .ip3(n1373), .ip4(n1226), .op(
        out[13]) );
  nor2_1 U1517 ( .ip1(n1229), .ip2(n2024), .op(n2023) );
  nand2_1 U1518 ( .ip1(n2022), .ip2(n1438), .op(n1236) );
  nor2_1 U1519 ( .ip1(in1[14]), .ip2(in2[0]), .op(n1230) );
  not_ab_or_c_or_d U1520 ( .ip1(in2[0]), .ip2(n1580), .ip3(n1230), .ip4(n1058), 
        .op(n1231) );
  not_ab_or_c_or_d U1521 ( .ip1(n2106), .ip2(in1[13]), .ip3(n1232), .ip4(n1231), .op(n1792) );
  inv_1 U1522 ( .ip(n1792), .op(n1365) );
  or2_1 U1523 ( .ip1(n1365), .ip2(n2024), .op(n1235) );
  nand2_1 U1524 ( .ip1(in2[3]), .ip2(n1233), .op(n1234) );
  and4_1 U1525 ( .ip1(n1893), .ip2(n1236), .ip3(n1235), .ip4(n1234), .op(n1241) );
  nor2_1 U1526 ( .ip1(n1131), .ip2(n1458), .op(n1239) );
  nor2_1 U1527 ( .ip1(n1237), .ip2(n2024), .op(n1238) );
  not_ab_or_c_or_d U1528 ( .ip1(n2022), .ip2(n1350), .ip3(n1239), .ip4(n1238), 
        .op(n2042) );
  nor2_1 U1529 ( .ip1(n2042), .ip2(n1907), .op(n1240) );
  not_ab_or_c_or_d U1530 ( .ip1(n1874), .ip2(n2023), .ip3(n1241), .ip4(n1240), 
        .op(n1255) );
  inv_1 U1531 ( .ip(n1324), .op(n1248) );
  nor2_1 U1532 ( .ip1(in2[12]), .ip2(n1985), .op(n1242) );
  not_ab_or_c_or_d U1533 ( .ip1(n2092), .ip2(in2[12]), .ip3(n2099), .ip4(n1242), .op(n1243) );
  nor2_1 U1534 ( .ip1(n1243), .ip2(n1661), .op(n1247) );
  nor2_1 U1535 ( .ip1(n1985), .ip2(in1[12]), .op(n1244) );
  nor2_1 U1536 ( .ip1(n2099), .ip2(n1244), .op(n1245) );
  inv_1 U1537 ( .ip(in2[12]), .op(n1624) );
  nor2_1 U1538 ( .ip1(n1245), .ip2(n1624), .op(n1246) );
  not_ab_or_c_or_d U1539 ( .ip1(n1248), .ip2(n2028), .ip3(n1247), .ip4(n1246), 
        .op(n1254) );
  nor2_1 U1540 ( .ip1(n2014), .ip2(n2001), .op(n1902) );
  inv_1 U1541 ( .ip(n1902), .op(n1253) );
  fulladder U1542 ( .a(in1[12]), .b(n1250), .ci(n1249), .co(n1223), .s(n1251)
         );
  nand2_1 U1543 ( .ip1(n1251), .ip2(n2131), .op(n1252) );
  nand4_1 U1544 ( .ip1(n1255), .ip2(n1254), .ip3(n1253), .ip4(n1252), .op(
        out[12]) );
  nor2_1 U1545 ( .ip1(n1509), .ip2(n1256), .op(n1258) );
  nor3_1 U1546 ( .ip1(n1258), .ip2(in2[3]), .ip3(n1257), .op(n1997) );
  nand2_1 U1547 ( .ip1(n2014), .ip2(n1259), .op(n1263) );
  nand2_1 U1548 ( .ip1(n1509), .ip2(n1260), .op(n1262) );
  nand2_1 U1549 ( .ip1(in2[3]), .ip2(n1806), .op(n1261) );
  nand4_1 U1550 ( .ip1(n2003), .ip2(n1263), .ip3(n1262), .ip4(n1261), .op(
        n1979) );
  nor2_1 U1551 ( .ip1(n1979), .ip2(n1907), .op(n1264) );
  inv_1 U1552 ( .ip(n1373), .op(n1387) );
  not_ab_or_c_or_d U1553 ( .ip1(n1874), .ip2(n1997), .ip3(n1264), .ip4(n1387), 
        .op(n1288) );
  inv_1 U1554 ( .ip(n1265), .op(n1983) );
  nor2_1 U1555 ( .ip1(n1983), .ip2(n1324), .op(n1271) );
  nor2_1 U1556 ( .ip1(in2[11]), .ip2(in1[11]), .op(n1266) );
  nor2_1 U1557 ( .ip1(n1266), .ip2(n2046), .op(n1270) );
  nor2_1 U1558 ( .ip1(in2[11]), .ip2(n1359), .op(n1658) );
  nand2_1 U1559 ( .ip1(in2[11]), .ip2(n1359), .op(n1659) );
  inv_1 U1560 ( .ip(n1659), .op(n1653) );
  nor2_1 U1561 ( .ip1(n1658), .ip2(n1653), .op(n1729) );
  nor2_1 U1562 ( .ip1(n1729), .ip2(n1985), .op(n1269) );
  inv_1 U1563 ( .ip(in2[11]), .op(n1267) );
  nor3_1 U1564 ( .ip1(n1989), .ip2(n1267), .ip3(n1359), .op(n1268) );
  nor4_1 U1565 ( .ip1(n1271), .ip2(n1270), .ip3(n1269), .ip4(n1268), .op(n1287) );
  fulladder U1566 ( .a(in1[11]), .b(n1273), .ci(n1272), .co(n1249), .s(n1274)
         );
  nand2_1 U1567 ( .ip1(n1274), .ip2(n2131), .op(n1286) );
  nor2_1 U1568 ( .ip1(n2003), .ip2(n1275), .op(n1281) );
  nor2_1 U1569 ( .ip1(n1661), .ip2(n2007), .op(n1276) );
  not_ab_or_c_or_d U1570 ( .ip1(n2048), .ip2(in1[11]), .ip3(n1277), .ip4(n1276), .op(n1279) );
  nand2_1 U1571 ( .ip1(n1279), .ip2(n1278), .op(n1814) );
  nor2_1 U1572 ( .ip1(n1814), .ip2(n2024), .op(n1280) );
  nor2_1 U1573 ( .ip1(n1281), .ip2(n1280), .op(n1284) );
  nand2_1 U1574 ( .ip1(n1394), .ip2(n2015), .op(n1283) );
  nand2_1 U1575 ( .ip1(n2022), .ip2(n1813), .op(n1282) );
  nand4_1 U1576 ( .ip1(n1284), .ip2(n1893), .ip3(n1283), .ip4(n1282), .op(
        n1285) );
  nand4_1 U1577 ( .ip1(n1288), .ip2(n1287), .ip3(n1286), .ip4(n1285), .op(
        out[11]) );
  or2_1 U1578 ( .ip1(in2[10]), .ip2(in1[10]), .op(n1292) );
  inv_1 U1579 ( .ip(in2[10]), .op(n1289) );
  nor2_1 U1580 ( .ip1(in1[10]), .ip2(n1289), .op(n1654) );
  nor2_1 U1581 ( .ip1(in2[10]), .ip2(n1391), .op(n1660) );
  nor2_1 U1582 ( .ip1(n1654), .ip2(n1660), .op(n1728) );
  nor2_1 U1583 ( .ip1(n1728), .ip2(n1985), .op(n1291) );
  nor3_1 U1584 ( .ip1(n1989), .ip2(n1391), .ip3(n1289), .op(n1290) );
  not_ab_or_c_or_d U1585 ( .ip1(n2099), .ip2(n1292), .ip3(n1291), .ip4(n1290), 
        .op(n1321) );
  fulladder U1586 ( .a(in1[10]), .b(n1294), .ci(n1293), .co(n1272), .s(n1316)
         );
  nor2_1 U1587 ( .ip1(n1295), .ip2(n1907), .op(n1315) );
  nor2_1 U1588 ( .ip1(n1468), .ip2(n2003), .op(n1313) );
  nand2_1 U1589 ( .ip1(n1297), .ip2(n1296), .op(n1300) );
  nand2_1 U1590 ( .ip1(n1298), .ip2(n1937), .op(n1299) );
  nand2_1 U1591 ( .ip1(n1300), .ip2(n1299), .op(n1466) );
  inv_1 U1592 ( .ip(n1466), .op(n1888) );
  nor2_1 U1593 ( .ip1(n1815), .ip2(n1888), .op(n1312) );
  nor2_1 U1594 ( .ip1(n1661), .ip2(n2102), .op(n1302) );
  nor2_1 U1595 ( .ip1(n1783), .ip2(n1554), .op(n1301) );
  nor4_1 U1596 ( .ip1(n1304), .ip2(n1303), .ip3(n1302), .ip4(n1301), .op(n1492) );
  nand2_1 U1597 ( .ip1(n2014), .ip2(n1492), .op(n1310) );
  nor2_1 U1598 ( .ip1(n1543), .ip2(n2102), .op(n1308) );
  nor2_1 U1599 ( .ip1(in1[15]), .ip2(in2[1]), .op(n1305) );
  not_ab_or_c_or_d U1600 ( .ip1(in2[1]), .ip2(n1306), .ip3(n1305), .ip4(n1772), 
        .op(n1307) );
  not_ab_or_c_or_d U1601 ( .ip1(n2048), .ip2(in1[14]), .ip3(n1308), .ip4(n1307), .op(n1891) );
  nand2_1 U1602 ( .ip1(n1891), .ip2(n2022), .op(n1309) );
  nand2_1 U1603 ( .ip1(n1310), .ip2(n1309), .op(n1311) );
  nor4_1 U1604 ( .ip1(n1313), .ip2(n1312), .ip3(n1854), .ip4(n1311), .op(n1314) );
  not_ab_or_c_or_d U1605 ( .ip1(n1316), .ip2(n2131), .ip3(n1315), .ip4(n1314), 
        .op(n1320) );
  nand2_1 U1606 ( .ip1(n1874), .ip2(n1317), .op(n1319) );
  or2_1 U1607 ( .ip1(n1324), .ip2(n1469), .op(n1318) );
  nand4_1 U1608 ( .ip1(n1321), .ip2(n1320), .ip3(n1319), .ip4(n1318), .op(
        out[10]) );
  inv_1 U1609 ( .ip(n1522), .op(n1332) );
  nor2_1 U1610 ( .ip1(n1322), .ip2(n1907), .op(n1331) );
  nor2_1 U1611 ( .ip1(in2[9]), .ip2(in1[9]), .op(n1323) );
  nor2_1 U1612 ( .ip1(n1323), .ip2(n2046), .op(n1329) );
  nand2_1 U1613 ( .ip1(in2[9]), .ip2(n1389), .op(n1652) );
  inv_1 U1614 ( .ip(in2[9]), .op(n1325) );
  nand2_1 U1615 ( .ip1(in1[9]), .ip2(n1325), .op(n1569) );
  and2_1 U1616 ( .ip1(n1652), .ip2(n1569), .op(n1727) );
  nor2_1 U1617 ( .ip1(n1727), .ip2(n1985), .op(n1328) );
  nor2_1 U1618 ( .ip1(n1521), .ip2(n1324), .op(n1327) );
  nor3_1 U1619 ( .ip1(n1989), .ip2(n1389), .ip3(n1325), .op(n1326) );
  or4_1 U1620 ( .ip1(n1329), .ip2(n1328), .ip3(n1327), .ip4(n1326), .op(n1330)
         );
  not_ab_or_c_or_d U1621 ( .ip1(n1845), .ip2(n1332), .ip3(n1331), .ip4(n1330), 
        .op(n1346) );
  nor2_1 U1622 ( .ip1(n1131), .ip2(n1333), .op(n1339) );
  nand2_1 U1623 ( .ip1(in1[11]), .ip2(n1508), .op(n1336) );
  nand2_1 U1624 ( .ip1(in1[9]), .ip2(n2048), .op(n1335) );
  nand2_1 U1625 ( .ip1(in1[10]), .ip2(n2106), .op(n1334) );
  nand4_1 U1626 ( .ip1(n1337), .ip2(n1336), .ip3(n1335), .ip4(n1334), .op(
        n1848) );
  nor2_1 U1627 ( .ip1(n1848), .ip2(n2024), .op(n1338) );
  not_ab_or_c_or_d U1628 ( .ip1(n2022), .ip2(n1852), .ip3(n1339), .ip4(n1338), 
        .op(n1340) );
  nand2_1 U1629 ( .ip1(n1893), .ip2(n1340), .op(n1345) );
  fulladder U1630 ( .a(in1[9]), .b(n1342), .ci(n1341), .co(n1293), .s(n1343)
         );
  nand2_1 U1631 ( .ip1(n1343), .ip2(n2131), .op(n1344) );
  nand4_1 U1632 ( .ip1(n1346), .ip2(n1373), .ip3(n1345), .ip4(n1344), .op(
        out[9]) );
  nor2_1 U1633 ( .ip1(n1131), .ip2(n1769), .op(n1349) );
  nor2_1 U1634 ( .ip1(n1347), .ip2(n1941), .op(n1348) );
  not_ab_or_c_or_d U1635 ( .ip1(n1350), .ip2(n2014), .ip3(n1349), .ip4(n1348), 
        .op(n1947) );
  nor2_1 U1636 ( .ip1(n1947), .ip2(n1907), .op(n1355) );
  nor2_1 U1637 ( .ip1(in2[8]), .ip2(in1[8]), .op(n1351) );
  nor2_1 U1638 ( .ip1(n1351), .ip2(n2046), .op(n1354) );
  xor2_1 U1639 ( .ip1(in2[8]), .ip2(n1567), .op(n1726) );
  nor2_1 U1640 ( .ip1(n1985), .ip2(n1726), .op(n1353) );
  inv_1 U1641 ( .ip(in2[8]), .op(n1564) );
  nor3_1 U1642 ( .ip1(n1989), .ip2(n1567), .ip3(n1564), .op(n1352) );
  nor4_1 U1643 ( .ip1(n1355), .ip2(n1354), .ip3(n1353), .ip4(n1352), .op(n1374) );
  fulladder U1644 ( .a(in1[8]), .b(n1357), .ci(n1356), .co(n1341), .s(n1358)
         );
  nand2_1 U1645 ( .ip1(n1358), .ip2(n2131), .op(n1372) );
  nor2_1 U1646 ( .ip1(n1359), .ip2(n1783), .op(n1360) );
  nor4_1 U1647 ( .ip1(n1363), .ip2(n1362), .ip3(n1361), .ip4(n1360), .op(n1789) );
  nor2_1 U1648 ( .ip1(n1789), .ip2(n1509), .op(n1364) );
  not_ab_or_c_or_d U1649 ( .ip1(in2[2]), .ip2(n1365), .ip3(in2[3]), .ip4(n1364), .op(n1366) );
  not_ab_or_c_or_d U1650 ( .ip1(in2[3]), .ip2(n1793), .ip3(in2[4]), .ip4(n1366), .op(n1369) );
  inv_1 U1651 ( .ip(n1962), .op(n1367) );
  nor3_1 U1652 ( .ip1(in2[3]), .ip2(n2100), .ip3(n1367), .op(n1368) );
  or2_1 U1653 ( .ip1(n1369), .ip2(n1368), .op(n1370) );
  nand2_1 U1654 ( .ip1(n1798), .ip2(n1370), .op(n1371) );
  nand4_1 U1655 ( .ip1(n1374), .ip2(n1373), .ip3(n1372), .ip4(n1371), .op(
        out[8]) );
  nor2_1 U1656 ( .ip1(in2[7]), .ip2(in1[7]), .op(n1375) );
  nor2_1 U1657 ( .ip1(n1375), .ip2(n2046), .op(n1380) );
  nand2_1 U1658 ( .ip1(in2[7]), .ip2(n1376), .op(n1647) );
  nor2_1 U1659 ( .ip1(in2[7]), .ip2(n1376), .op(n1646) );
  inv_1 U1660 ( .ip(n1646), .op(n1563) );
  nand2_1 U1661 ( .ip1(n1647), .ip2(n1563), .op(n1746) );
  nand2_1 U1662 ( .ip1(n2096), .ip2(n1746), .op(n1378) );
  nand3_1 U1663 ( .ip1(n2092), .ip2(in2[7]), .ip3(in1[7]), .op(n1377) );
  nand2_1 U1664 ( .ip1(n1378), .ip2(n1377), .op(n1379) );
  not_ab_or_c_or_d U1665 ( .ip1(n1876), .ip2(n1381), .ip3(n1380), .ip4(n1379), 
        .op(n1405) );
  fulladder U1666 ( .a(in1[7]), .b(n1383), .ci(n1382), .co(n1356), .s(n1388)
         );
  nand2_1 U1667 ( .ip1(n2124), .ip2(n1384), .op(n1840) );
  nor2_1 U1668 ( .ip1(n1840), .ip2(n1385), .op(n1386) );
  not_ab_or_c_or_d U1669 ( .ip1(n1388), .ip2(n2131), .ip3(n1387), .ip4(n1386), 
        .op(n1404) );
  nor2_1 U1670 ( .ip1(n1389), .ip2(n2102), .op(n1393) );
  nor2_1 U1671 ( .ip1(in1[8]), .ip2(in2[1]), .op(n1390) );
  not_ab_or_c_or_d U1672 ( .ip1(in2[1]), .ip2(n1391), .ip3(n1390), .ip4(n1772), 
        .op(n1392) );
  not_ab_or_c_or_d U1673 ( .ip1(n2048), .ip2(in1[7]), .ip3(n1393), .ip4(n1392), 
        .op(n1820) );
  nor2_1 U1674 ( .ip1(n1941), .ip2(n1814), .op(n1398) );
  nand2_1 U1675 ( .ip1(n1813), .ip2(n2015), .op(n1396) );
  nand2_1 U1676 ( .ip1(n1394), .ip2(n1946), .op(n1395) );
  nand2_1 U1677 ( .ip1(n1396), .ip2(n1395), .op(n1397) );
  not_ab_or_c_or_d U1678 ( .ip1(n2014), .ip2(n1820), .ip3(n1398), .ip4(n1397), 
        .op(n1399) );
  nand2_1 U1679 ( .ip1(n1893), .ip2(n1399), .op(n1403) );
  inv_1 U1680 ( .ip(n1400), .op(n1401) );
  nand2_1 U1681 ( .ip1(n1845), .ip2(n1401), .op(n1402) );
  nand4_1 U1682 ( .ip1(n1405), .ip2(n1404), .ip3(n1403), .ip4(n1402), .op(
        out[7]) );
  or2_1 U1683 ( .ip1(in2[6]), .ip2(in1[6]), .op(n1415) );
  nor2_1 U1684 ( .ip1(n1840), .ip2(n1406), .op(n1414) );
  nor2_1 U1685 ( .ip1(in2[6]), .ip2(n1407), .op(n1648) );
  inv_1 U1686 ( .ip(in2[6]), .op(n1408) );
  nor2_1 U1687 ( .ip1(in1[6]), .ip2(n1408), .op(n1643) );
  or2_1 U1688 ( .ip1(n1648), .ip2(n1643), .op(n1745) );
  nand2_1 U1689 ( .ip1(n2096), .ip2(n1745), .op(n1412) );
  nand2_1 U1690 ( .ip1(n1876), .ip2(n1409), .op(n1411) );
  nand3_1 U1691 ( .ip1(n2092), .ip2(in1[6]), .ip3(in2[6]), .op(n1410) );
  nand3_1 U1692 ( .ip1(n1412), .ip2(n1411), .ip3(n1410), .op(n1413) );
  not_ab_or_c_or_d U1693 ( .ip1(n2099), .ip2(n1415), .ip3(n1414), .ip4(n1413), 
        .op(n1432) );
  nand4_1 U1694 ( .ip1(n1419), .ip2(n1418), .ip3(n1417), .ip4(n1416), .op(
        n1489) );
  nor2_1 U1695 ( .ip1(n1489), .ip2(n2024), .op(n1423) );
  nand2_1 U1696 ( .ip1(n2022), .ip2(n1492), .op(n1421) );
  nand2_1 U1697 ( .ip1(n1891), .ip2(n2015), .op(n1420) );
  nand2_1 U1698 ( .ip1(n1421), .ip2(n1420), .op(n1422) );
  not_ab_or_c_or_d U1699 ( .ip1(n1466), .ip2(n1946), .ip3(n1423), .ip4(n1422), 
        .op(n1424) );
  nand2_1 U1700 ( .ip1(n1893), .ip2(n1424), .op(n1431) );
  fulladder U1701 ( .a(in1[6]), .b(n1426), .ci(n1425), .co(n1382), .s(n1427)
         );
  nand2_1 U1702 ( .ip1(n1427), .ip2(n2131), .op(n1430) );
  inv_1 U1703 ( .ip(n1874), .op(n1843) );
  or2_1 U1704 ( .ip1(n1428), .ip2(n1843), .op(n1429) );
  nand4_1 U1705 ( .ip1(n1432), .ip2(n1431), .ip3(n1430), .ip4(n1429), .op(
        out[6]) );
  nor2_1 U1706 ( .ip1(n1807), .ip2(n1989), .op(n1437) );
  nor2_1 U1707 ( .ip1(in2[4]), .ip2(in1[4]), .op(n1433) );
  nor2_1 U1708 ( .ip1(n1433), .ip2(n2046), .op(n1436) );
  nor2_1 U1709 ( .ip1(in2[4]), .ip2(n1807), .op(n1641) );
  nor2_1 U1710 ( .ip1(in1[4]), .ip2(n2100), .op(n1637) );
  or2_1 U1711 ( .ip1(n1641), .ip2(n1637), .op(n1704) );
  inv_1 U1712 ( .ip(n1704), .op(n1434) );
  nor2_1 U1713 ( .ip1(n1434), .ip2(n1985), .op(n1435) );
  not_ab_or_c_or_d U1714 ( .ip1(in2[4]), .ip2(n1437), .ip3(n1436), .ip4(n1435), 
        .op(n1462) );
  nand2_1 U1715 ( .ip1(n1438), .ip2(n1946), .op(n1445) );
  nand2_1 U1716 ( .ip1(n1789), .ip2(n2022), .op(n1444) );
  nor4_1 U1717 ( .ip1(n1442), .ip2(n1441), .ip3(n1440), .ip4(n1439), .op(n1795) );
  nand2_1 U1718 ( .ip1(n1795), .ip2(n2014), .op(n1443) );
  nand3_1 U1719 ( .ip1(n1445), .ip2(n1444), .ip3(n1443), .op(n1446) );
  not_ab_or_c_or_d U1720 ( .ip1(n1792), .ip2(n2015), .ip3(n1446), .ip4(n1854), 
        .op(n1454) );
  nor2_1 U1721 ( .ip1(n1447), .ip2(n1843), .op(n1450) );
  nor2_1 U1722 ( .ip1(n1448), .ip2(n1821), .op(n1449) );
  nor2_1 U1723 ( .ip1(n1450), .ip2(n1449), .op(n1451) );
  nor2_1 U1724 ( .ip1(n1452), .ip2(n1451), .op(n1453) );
  nor2_1 U1725 ( .ip1(n1454), .ip2(n1453), .op(n1461) );
  fulladder U1726 ( .a(in1[4]), .b(n1456), .ci(n1455), .co(n1862), .s(n1457)
         );
  nand2_1 U1727 ( .ip1(n1457), .ip2(n2131), .op(n1460) );
  or2_1 U1728 ( .ip1(n1458), .ip2(n1840), .op(n1459) );
  nand4_1 U1729 ( .ip1(n1462), .ip2(n1461), .ip3(n1460), .ip4(n1459), .op(
        out[4]) );
  fulladder U1730 ( .a(in1[2]), .b(n1464), .ci(n1463), .co(n1826), .s(n1477)
         );
  nor2_1 U1731 ( .ip1(n1509), .ip2(in1[2]), .op(n1465) );
  nor2_1 U1732 ( .ip1(n1465), .ip2(n2046), .op(n1476) );
  nor2_1 U1733 ( .ip1(n1509), .ip2(n1472), .op(n1635) );
  nor2_1 U1734 ( .ip1(in1[2]), .ip2(n1149), .op(n1630) );
  or2_1 U1735 ( .ip1(n1635), .ip2(n1630), .op(n1703) );
  nor2_1 U1736 ( .ip1(n1466), .ip2(n1509), .op(n1467) );
  not_ab_or_c_or_d U1737 ( .ip1(in2[2]), .ip2(n1468), .ip3(in2[3]), .ip4(n1467), .op(n1482) );
  inv_1 U1738 ( .ip(n1482), .op(n1471) );
  nand2_1 U1739 ( .ip1(in2[3]), .ip2(n1469), .op(n1470) );
  nand2_1 U1740 ( .ip1(n1471), .ip2(n1470), .op(n1913) );
  nor2_1 U1741 ( .ip1(n1913), .ip2(n1821), .op(n1474) );
  nor3_1 U1742 ( .ip1(n1989), .ip2(n1149), .ip3(n1472), .op(n1473) );
  ab_or_c_or_d U1743 ( .ip1(n2096), .ip2(n1703), .ip3(n1474), .ip4(n1473), 
        .op(n1475) );
  not_ab_or_c_or_d U1744 ( .ip1(n1477), .ip2(n2131), .ip3(n1476), .ip4(n1475), 
        .op(n1498) );
  nor2_1 U1745 ( .ip1(n1479), .ip2(n1478), .op(n1480) );
  nor2_1 U1746 ( .ip1(n1480), .ip2(n1131), .op(n1481) );
  nor2_1 U1747 ( .ip1(n1482), .ip2(n1481), .op(n1923) );
  nand2_1 U1748 ( .ip1(n1874), .ip2(n1923), .op(n1497) );
  nor2_1 U1749 ( .ip1(in2[2]), .ip2(n1840), .op(n1839) );
  inv_1 U1750 ( .ip(n1927), .op(n1483) );
  nand2_1 U1751 ( .ip1(n1839), .ip2(n1483), .op(n1496) );
  nor2_1 U1752 ( .ip1(in1[3]), .ip2(n2007), .op(n1485) );
  nor2_1 U1753 ( .ip1(in1[2]), .ip2(n1782), .op(n1484) );
  not_ab_or_c_or_d U1754 ( .ip1(n1486), .ip2(n1857), .ip3(n1485), .ip4(n1484), 
        .op(n1488) );
  nand2_1 U1755 ( .ip1(n1508), .ip2(n1807), .op(n1487) );
  not_ab_or_c_or_d U1756 ( .ip1(n1488), .ip2(n1487), .ip3(in2[3]), .ip4(n1509), 
        .op(n1491) );
  nor2_1 U1757 ( .ip1(n1941), .ip2(n1489), .op(n1490) );
  not_ab_or_c_or_d U1758 ( .ip1(n1492), .ip2(n2015), .ip3(n1491), .ip4(n1490), 
        .op(n1494) );
  nand2_1 U1759 ( .ip1(n1891), .ip2(n1946), .op(n1493) );
  nand3_1 U1760 ( .ip1(n1893), .ip2(n1494), .ip3(n1493), .op(n1495) );
  nand4_1 U1761 ( .ip1(n1498), .ip2(n1497), .ip3(n1496), .ip4(n1495), .op(
        out[2]) );
  nand2_1 U1762 ( .ip1(n1499), .ip2(n1058), .op(n1502) );
  nor2_1 U1763 ( .ip1(in1[1]), .ip2(n1058), .op(n1632) );
  nor2_1 U1764 ( .ip1(in2[1]), .ip2(n1499), .op(n1557) );
  nor2_1 U1765 ( .ip1(n1632), .ip2(n1557), .op(n1708) );
  nor2_1 U1766 ( .ip1(n1708), .ip2(n1985), .op(n1501) );
  nor3_1 U1767 ( .ip1(n1989), .ip2(n1499), .ip3(n1058), .op(n1500) );
  not_ab_or_c_or_d U1768 ( .ip1(n2099), .ip2(n1502), .ip3(n1501), .ip4(n1500), 
        .op(n1536) );
  nor2_1 U1769 ( .ip1(in1[6]), .ip2(in2[1]), .op(n1503) );
  not_ab_or_c_or_d U1770 ( .ip1(in2[1]), .ip2(n1567), .ip3(n1503), .ip4(n1772), 
        .op(n1504) );
  not_ab_or_c_or_d U1771 ( .ip1(n1508), .ip2(in1[7]), .ip3(n1505), .ip4(n1504), 
        .op(n1855) );
  inv_1 U1772 ( .ip(in1[3]), .op(n1830) );
  nor2_1 U1773 ( .ip1(in1[2]), .ip2(n2007), .op(n1507) );
  nor2_1 U1774 ( .ip1(in1[1]), .ip2(n1782), .op(n1506) );
  not_ab_or_c_or_d U1775 ( .ip1(n1508), .ip2(n1830), .ip3(n1507), .ip4(n1506), 
        .op(n1511) );
  not_ab_or_c_or_d U1776 ( .ip1(n1511), .ip2(n1510), .ip3(in2[3]), .ip4(n1509), 
        .op(n1514) );
  nor2_1 U1777 ( .ip1(n1852), .ip2(n1149), .op(n1512) );
  not_ab_or_c_or_d U1778 ( .ip1(n1848), .ip2(n1149), .ip3(n1131), .ip4(n1512), 
        .op(n1513) );
  not_ab_or_c_or_d U1779 ( .ip1(n2022), .ip2(n1855), .ip3(n1514), .ip4(n1513), 
        .op(n1515) );
  nor2_1 U1780 ( .ip1(in2[4]), .ip2(n1515), .op(n1520) );
  inv_1 U1781 ( .ip(n1798), .op(n1517) );
  nor2_1 U1782 ( .ip1(n1517), .ip2(n1516), .op(n1518) );
  nor2_1 U1783 ( .ip1(n1893), .ip2(n1518), .op(n1519) );
  nor2_1 U1784 ( .ip1(n1520), .ip2(n1519), .op(n1527) );
  nor2_1 U1785 ( .ip1(n1521), .ip2(n1821), .op(n1524) );
  nor2_1 U1786 ( .ip1(n1522), .ip2(n1843), .op(n1523) );
  nor2_1 U1787 ( .ip1(n1524), .ip2(n1523), .op(n1525) );
  nor2_1 U1788 ( .ip1(n1525), .ip2(n1131), .op(n1526) );
  nor2_1 U1789 ( .ip1(n1527), .ip2(n1526), .op(n1535) );
  inv_1 U1790 ( .ip(n1528), .op(n1529) );
  nand2_1 U1791 ( .ip1(n1529), .ip2(n1839), .op(n1534) );
  fulladder U1792 ( .a(in1[1]), .b(n1531), .ci(n1530), .co(n1463), .s(n1532)
         );
  nand2_1 U1793 ( .ip1(n1532), .ip2(n2131), .op(n1533) );
  nand4_1 U1794 ( .ip1(n1536), .ip2(n1535), .ip3(n1534), .ip4(n1533), .op(
        out[1]) );
  inv_1 U1795 ( .ip(in2[31]), .op(n1537) );
  nor2_1 U1796 ( .ip1(N316), .ip2(n1537), .op(n1760) );
  inv_1 U1797 ( .ip(in1[28]), .op(n1538) );
  nor2_1 U1798 ( .ip1(in2[28]), .ip2(n1538), .op(n1713) );
  nor2_1 U1799 ( .ip1(in2[29]), .ip2(n2103), .op(n1690) );
  inv_1 U1800 ( .ip(n1690), .op(n1711) );
  nand2_1 U1801 ( .ip1(n1539), .ip2(n1711), .op(n1540) );
  nor2_1 U1802 ( .ip1(n1713), .ip2(n1540), .op(n1592) );
  inv_1 U1803 ( .ip(in2[27]), .op(n1988) );
  nor2_1 U1804 ( .ip1(in1[27]), .ip2(n1988), .op(n1720) );
  nand2_1 U1805 ( .ip1(in2[24]), .ip2(n1952), .op(n1681) );
  inv_1 U1806 ( .ip(n1681), .op(n1722) );
  inv_1 U1807 ( .ip(n1602), .op(n1542) );
  not_ab_or_c_or_d U1808 ( .ip1(n1722), .ip2(n1542), .ip3(n1541), .ip4(n1683), 
        .op(n1589) );
  inv_1 U1809 ( .ip(n1617), .op(n1551) );
  nor2_1 U1810 ( .ip1(n1613), .ip2(n1610), .op(n1669) );
  inv_1 U1811 ( .ip(in2[18]), .op(n1914) );
  nor2_1 U1812 ( .ip1(in1[18]), .ip2(n1914), .op(n1731) );
  inv_1 U1813 ( .ip(n1606), .op(n1546) );
  nand3_1 U1814 ( .ip1(in2[16]), .ip2(n1543), .ip3(n1605), .op(n1544) );
  nor2_1 U1815 ( .ip1(in2[18]), .ip2(n1915), .op(n1730) );
  not_ab_or_c_or_d U1816 ( .ip1(n1674), .ip2(n1544), .ip3(n1730), .ip4(n1606), 
        .op(n1545) );
  not_ab_or_c_or_d U1817 ( .ip1(n1731), .ip2(n1546), .ip3(n1620), .ip4(n1545), 
        .op(n1547) );
  or2_1 U1818 ( .ip1(n1552), .ip2(n1547), .op(n1549) );
  nor2_1 U1819 ( .ip1(n1617), .ip2(n1619), .op(n1584) );
  inv_1 U1820 ( .ip(n1584), .op(n1548) );
  not_ab_or_c_or_d U1821 ( .ip1(n1669), .ip2(n1549), .ip3(n1553), .ip4(n1548), 
        .op(n1550) );
  not_ab_or_c_or_d U1822 ( .ip1(n1611), .ip2(n1551), .ip3(n1550), .ip4(n1612), 
        .op(n1587) );
  nor2_1 U1823 ( .ip1(n1553), .ip2(n1552), .op(n1615) );
  nor2_1 U1824 ( .ip1(n1606), .ip2(n1730), .op(n1585) );
  inv_1 U1825 ( .ip(in2[14]), .op(n1880) );
  nor2_1 U1826 ( .ip1(n1880), .ip2(in1[14]), .op(n1621) );
  nand2_1 U1827 ( .ip1(in2[13]), .ip2(n1554), .op(n1663) );
  nand3_1 U1828 ( .ip1(in2[12]), .ip2(n1661), .ip3(n1623), .op(n1555) );
  nor2_1 U1829 ( .ip1(in2[14]), .ip2(n1882), .op(n1885) );
  not_ab_or_c_or_d U1830 ( .ip1(n1663), .ip2(n1555), .ip3(n1574), .ip4(n1885), 
        .op(n1579) );
  inv_1 U1831 ( .ip(n1658), .op(n1573) );
  nor2_1 U1832 ( .ip1(in2[5]), .ip2(n1857), .op(n1640) );
  inv_1 U1833 ( .ip(n1640), .op(n1699) );
  nor2_1 U1834 ( .ip1(in2[3]), .ip2(n1830), .op(n1634) );
  inv_1 U1835 ( .ip(n1634), .op(n1701) );
  inv_1 U1836 ( .ip(n1706), .op(n1775) );
  nor2_1 U1837 ( .ip1(n1632), .ip2(n1775), .op(n1556) );
  nor4_1 U1838 ( .ip1(n1634), .ip2(n1635), .ip3(n1557), .ip4(n1556), .op(n1558) );
  nand2_1 U1839 ( .ip1(in2[3]), .ip2(n1830), .op(n1702) );
  inv_1 U1840 ( .ip(n1702), .op(n1631) );
  not_ab_or_c_or_d U1841 ( .ip1(n1630), .ip2(n1701), .ip3(n1558), .ip4(n1631), 
        .op(n1559) );
  nor3_1 U1842 ( .ip1(n1640), .ip2(n1641), .ip3(n1559), .op(n1560) );
  nand2_1 U1843 ( .ip1(in2[5]), .ip2(n1857), .op(n1700) );
  inv_1 U1844 ( .ip(n1700), .op(n1638) );
  not_ab_or_c_or_d U1845 ( .ip1(n1637), .ip2(n1699), .ip3(n1560), .ip4(n1638), 
        .op(n1561) );
  nor3_1 U1846 ( .ip1(n1646), .ip2(n1648), .ip3(n1561), .op(n1562) );
  inv_1 U1847 ( .ip(n1647), .op(n1644) );
  not_ab_or_c_or_d U1848 ( .ip1(n1643), .ip2(n1563), .ip3(n1562), .ip4(n1644), 
        .op(n1566) );
  nand2_1 U1849 ( .ip1(in1[8]), .ip2(n1564), .op(n1565) );
  nand2_1 U1850 ( .ip1(n1569), .ip2(n1565), .op(n1651) );
  or2_1 U1851 ( .ip1(n1566), .ip2(n1651), .op(n1571) );
  nand2_1 U1852 ( .ip1(in2[8]), .ip2(n1567), .op(n1568) );
  nand2_1 U1853 ( .ip1(n1652), .ip2(n1568), .op(n1649) );
  nand2_1 U1854 ( .ip1(n1649), .ip2(n1569), .op(n1570) );
  not_ab_or_c_or_d U1855 ( .ip1(n1571), .ip2(n1570), .ip3(n1660), .ip4(n1658), 
        .op(n1572) );
  not_ab_or_c_or_d U1856 ( .ip1(n1654), .ip2(n1573), .ip3(n1653), .ip4(n1572), 
        .op(n1577) );
  nor2_1 U1857 ( .ip1(n1574), .ip2(n1885), .op(n1576) );
  nand2_1 U1858 ( .ip1(in1[12]), .ip2(n1624), .op(n1575) );
  nand3_1 U1859 ( .ip1(n1576), .ip2(n1623), .ip3(n1575), .op(n1710) );
  nor2_1 U1860 ( .ip1(n1577), .ip2(n1710), .op(n1578) );
  not_ab_or_c_or_d U1861 ( .ip1(n1621), .ip2(n1672), .ip3(n1579), .ip4(n1578), 
        .op(n1582) );
  nand2_1 U1862 ( .ip1(in2[15]), .ip2(n1580), .op(n1668) );
  inv_1 U1863 ( .ip(n1605), .op(n1581) );
  not_ab_or_c_or_d U1864 ( .ip1(n1582), .ip2(n1668), .ip3(n1603), .ip4(n1581), 
        .op(n1583) );
  nand4_1 U1865 ( .ip1(n1615), .ip2(n1585), .ip3(n1584), .ip4(n1583), .op(
        n1586) );
  nor2_1 U1866 ( .ip1(in2[24]), .ip2(n1952), .op(n1723) );
  ab_or_c_or_d U1867 ( .ip1(n1587), .ip2(n1586), .ip3(n1602), .ip4(n1723), 
        .op(n1588) );
  inv_1 U1868 ( .ip(in1[27]), .op(n1987) );
  nor2_1 U1869 ( .ip1(in2[27]), .ip2(n1987), .op(n1721) );
  not_ab_or_c_or_d U1870 ( .ip1(n1589), .ip2(n1588), .ip3(n1601), .ip4(n1721), 
        .op(n1590) );
  or2_1 U1871 ( .ip1(n1720), .ip2(n1590), .op(n1591) );
  nand2_1 U1872 ( .ip1(n1592), .ip2(n1591), .op(n1749) );
  nor2_1 U1873 ( .ip1(in2[31]), .ip2(n2093), .op(n1755) );
  or2_1 U1874 ( .ip1(n1749), .ip2(n1755), .op(n1597) );
  inv_1 U1875 ( .ip(in2[28]), .op(n1593) );
  nor2_1 U1876 ( .ip1(in1[28]), .ip2(n1593), .op(n1714) );
  nand2_1 U1877 ( .ip1(in2[29]), .ip2(n2103), .op(n1712) );
  inv_1 U1878 ( .ip(n1712), .op(n1594) );
  inv_1 U1879 ( .ip(n1599), .op(n1692) );
  not_ab_or_c_or_d U1880 ( .ip1(n1714), .ip2(n1711), .ip3(n1594), .ip4(n1692), 
        .op(n1595) );
  or2_1 U1881 ( .ip1(n1689), .ip2(n1595), .op(n1750) );
  or2_1 U1882 ( .ip1(n1750), .ip2(n1755), .op(n1596) );
  nand2_1 U1883 ( .ip1(n1597), .ip2(n1596), .op(n1598) );
  nor3_1 U1884 ( .ip1(op[0]), .ip2(n1760), .ip3(n1598), .op(n1698) );
  nand2_1 U1885 ( .ip1(n1599), .ip2(n1712), .op(n1600) );
  nor2_1 U1886 ( .ip1(n1714), .ip2(n1600), .op(n1688) );
  not_ab_or_c_or_d U1887 ( .ip1(n1723), .ip2(n1682), .ip3(n1602), .ip4(n1601), 
        .op(n1685) );
  nand2_1 U1888 ( .ip1(n1603), .ip2(n1674), .op(n1604) );
  not_ab_or_c_or_d U1889 ( .ip1(n1605), .ip2(n1604), .ip3(n1620), .ip4(n1731), 
        .op(n1607) );
  not_ab_or_c_or_d U1890 ( .ip1(n1730), .ip2(n1608), .ip3(n1607), .ip4(n1606), 
        .op(n1609) );
  or2_1 U1891 ( .ip1(n1610), .ip2(n1609), .op(n1614) );
  or2_1 U1892 ( .ip1(n1612), .ip2(n1611), .op(n1671) );
  not_ab_or_c_or_d U1893 ( .ip1(n1615), .ip2(n1614), .ip3(n1613), .ip4(n1671), 
        .op(n1616) );
  not_ab_or_c_or_d U1894 ( .ip1(n1619), .ip2(n1618), .ip3(n1617), .ip4(n1616), 
        .op(n1679) );
  nor2_1 U1895 ( .ip1(n1620), .ip2(n1731), .op(n1677) );
  inv_1 U1896 ( .ip(n1668), .op(n1622) );
  nor2_1 U1897 ( .ip1(n1622), .ip2(n1621), .op(n1664) );
  inv_1 U1898 ( .ip(n1664), .op(n1625) );
  or2_1 U1899 ( .ip1(n1623), .ip2(n1625), .op(n1628) );
  nand3_1 U1900 ( .ip1(in1[12]), .ip2(n1663), .ip3(n1624), .op(n1626) );
  or2_1 U1901 ( .ip1(n1626), .ip2(n1625), .op(n1627) );
  nand2_1 U1902 ( .ip1(n1628), .ip2(n1627), .op(n1667) );
  not_ab_or_c_or_d U1903 ( .ip1(in1[1]), .ip2(n1058), .ip3(in1[0]), .ip4(n1772), .op(n1629) );
  nor4_1 U1904 ( .ip1(n1632), .ip2(n1631), .ip3(n1630), .ip4(n1629), .op(n1633) );
  not_ab_or_c_or_d U1905 ( .ip1(n1635), .ip2(n1702), .ip3(n1634), .ip4(n1633), 
        .op(n1636) );
  nor3_1 U1906 ( .ip1(n1638), .ip2(n1637), .ip3(n1636), .op(n1639) );
  not_ab_or_c_or_d U1907 ( .ip1(n1641), .ip2(n1700), .ip3(n1640), .ip4(n1639), 
        .op(n1642) );
  nor3_1 U1908 ( .ip1(n1644), .ip2(n1643), .ip3(n1642), .op(n1645) );
  not_ab_or_c_or_d U1909 ( .ip1(n1648), .ip2(n1647), .ip3(n1646), .ip4(n1645), 
        .op(n1650) );
  or2_1 U1910 ( .ip1(n1650), .ip2(n1649), .op(n1656) );
  nand2_1 U1911 ( .ip1(n1652), .ip2(n1651), .op(n1655) );
  not_ab_or_c_or_d U1912 ( .ip1(n1656), .ip2(n1655), .ip3(n1654), .ip4(n1653), 
        .op(n1657) );
  not_ab_or_c_or_d U1913 ( .ip1(n1660), .ip2(n1659), .ip3(n1658), .ip4(n1657), 
        .op(n1665) );
  nand2_1 U1914 ( .ip1(in2[12]), .ip2(n1661), .op(n1662) );
  nand3_1 U1915 ( .ip1(n1664), .ip2(n1663), .ip3(n1662), .op(n1709) );
  nor2_1 U1916 ( .ip1(n1665), .ip2(n1709), .op(n1666) );
  not_ab_or_c_or_d U1917 ( .ip1(n1885), .ip2(n1668), .ip3(n1667), .ip4(n1666), 
        .op(n1673) );
  inv_1 U1918 ( .ip(n1669), .op(n1670) );
  not_ab_or_c_or_d U1919 ( .ip1(n1673), .ip2(n1672), .ip3(n1671), .ip4(n1670), 
        .op(n1676) );
  nand4_1 U1920 ( .ip1(n1677), .ip2(n1676), .ip3(n1675), .ip4(n1674), .op(
        n1678) );
  nand2_1 U1921 ( .ip1(n1679), .ip2(n1678), .op(n1680) );
  nand3_1 U1922 ( .ip1(n1682), .ip2(n1681), .ip3(n1680), .op(n1684) );
  not_ab_or_c_or_d U1923 ( .ip1(n1685), .ip2(n1684), .ip3(n1683), .ip4(n1720), 
        .op(n1686) );
  or2_1 U1924 ( .ip1(n1721), .ip2(n1686), .op(n1687) );
  nand2_1 U1925 ( .ip1(n1688), .ip2(n1687), .op(n1754) );
  or2_1 U1926 ( .ip1(n1754), .ip2(n1760), .op(n1694) );
  not_ab_or_c_or_d U1927 ( .ip1(n1713), .ip2(n1712), .ip3(n1690), .ip4(n1689), 
        .op(n1691) );
  or2_1 U1928 ( .ip1(n1692), .ip2(n1691), .op(n1756) );
  or2_1 U1929 ( .ip1(n1756), .ip2(n1760), .op(n1693) );
  nand2_1 U1930 ( .ip1(n1694), .ip2(n1693), .op(n1695) );
  nor3_1 U1931 ( .ip1(n1755), .ip2(n1748), .ip3(n1695), .op(n1697) );
  or4_1 U1932 ( .ip1(n1698), .ip2(n1697), .ip3(n1696), .ip4(n1771), .op(n1768)
         );
  nand2_1 U1933 ( .ip1(n1700), .ip2(n1699), .op(n1861) );
  nand2_1 U1934 ( .ip1(n1702), .ip2(n1701), .op(n1825) );
  nor4_1 U1935 ( .ip1(n1861), .ip2(n1704), .ip3(n1825), .ip4(n1703), .op(n1707) );
  nand2_1 U1936 ( .ip1(in1[0]), .ip2(n1772), .op(n1705) );
  nand4_1 U1937 ( .ip1(n1708), .ip2(n1707), .ip3(n1706), .ip4(n1705), .op(
        n1744) );
  inv_1 U1938 ( .ip(n1709), .op(n1742) );
  inv_1 U1939 ( .ip(n1710), .op(n1741) );
  or2_1 U1940 ( .ip1(n1755), .ip2(n1760), .op(n2095) );
  nand2_1 U1941 ( .ip1(n1712), .ip2(n1711), .op(n2067) );
  or2_1 U1942 ( .ip1(n1714), .ip2(n1713), .op(n2026) );
  nor4_1 U1943 ( .ip1(n2095), .ip2(n1715), .ip3(n2067), .ip4(n2026), .op(n1740) );
  nand4_1 U1944 ( .ip1(n1719), .ip2(n1718), .ip3(n1717), .ip4(n1716), .op(
        n1738) );
  nor2_1 U1945 ( .ip1(n1721), .ip2(n1720), .op(n1986) );
  nor2_1 U1946 ( .ip1(n1723), .ip2(n1722), .op(n1951) );
  nand4_1 U1947 ( .ip1(n1986), .ip2(n1725), .ip3(n1724), .ip4(n1951), .op(
        n1737) );
  nand4_1 U1948 ( .ip1(n1729), .ip2(n1728), .ip3(n1727), .ip4(n1726), .op(
        n1736) );
  nor2_1 U1949 ( .ip1(n1731), .ip2(n1730), .op(n1911) );
  nand4_1 U1950 ( .ip1(n1734), .ip2(n1911), .ip3(n1733), .ip4(n1732), .op(
        n1735) );
  nor4_1 U1951 ( .ip1(n1738), .ip2(n1737), .ip3(n1736), .ip4(n1735), .op(n1739) );
  nand4_1 U1952 ( .ip1(n1742), .ip2(n1741), .ip3(n1740), .ip4(n1739), .op(
        n1743) );
  nor4_1 U1953 ( .ip1(n1746), .ip2(n1745), .ip3(n1744), .ip4(n1743), .op(n1747) );
  mux2_1 U1954 ( .ip1(op[0]), .ip2(n1748), .s(n1747), .op(n1765) );
  or2_1 U1955 ( .ip1(n1749), .ip2(n1760), .op(n1752) );
  or2_1 U1956 ( .ip1(n1750), .ip2(n1760), .op(n1751) );
  nand2_1 U1957 ( .ip1(n1752), .ip2(n1751), .op(n1753) );
  nor2_1 U1958 ( .ip1(n1755), .ip2(n1753), .op(n1762) );
  or2_1 U1959 ( .ip1(n1754), .ip2(n1755), .op(n1758) );
  or2_1 U1960 ( .ip1(n1756), .ip2(n1755), .op(n1757) );
  nand2_1 U1961 ( .ip1(n1758), .ip2(n1757), .op(n1759) );
  nor2_1 U1962 ( .ip1(n1760), .ip2(n1759), .op(n1761) );
  mux2_1 U1963 ( .ip1(n1762), .ip2(n1761), .s(op[0]), .op(n1763) );
  inv_1 U1964 ( .ip(n1763), .op(n1764) );
  mux2_1 U1965 ( .ip1(n1765), .ip2(n1764), .s(op[2]), .op(n1766) );
  nand2_1 U1966 ( .ip1(n1771), .ip2(n1766), .op(n1767) );
  nand2_1 U1967 ( .ip1(n1768), .ip2(n1767), .op(n1781) );
  nor2_1 U1968 ( .ip1(n1769), .ip2(n1840), .op(n1780) );
  nand2_1 U1969 ( .ip1(in2[0]), .ip2(n2099), .op(n1778) );
  not_ab_or_c_or_d U1970 ( .ip1(in2[0]), .ip2(n1771), .ip3(op[3]), .ip4(n1770), 
        .op(n1774) );
  nand2_1 U1971 ( .ip1(op[0]), .ip2(n1772), .op(n1773) );
  nand3_1 U1972 ( .ip1(op[2]), .ip2(n1774), .ip3(n1773), .op(n1777) );
  nand2_1 U1973 ( .ip1(n1775), .ip2(n2096), .op(n1776) );
  nand3_1 U1974 ( .ip1(n1778), .ip2(n1777), .ip3(n1776), .op(n1779) );
  not_ab_or_c_or_d U1975 ( .ip1(op[3]), .ip2(n1781), .ip3(n1780), .ip4(n1779), 
        .op(n1805) );
  nor2_1 U1976 ( .ip1(in1[2]), .ip2(n2102), .op(n1787) );
  nor2_1 U1977 ( .ip1(in1[0]), .ip2(n1782), .op(n1786) );
  nor2_1 U1978 ( .ip1(in1[3]), .ip2(n1783), .op(n1785) );
  nor2_1 U1979 ( .ip1(in1[1]), .ip2(n2007), .op(n1784) );
  nor4_1 U1980 ( .ip1(n1787), .ip2(n1786), .ip3(n1785), .ip4(n1784), .op(n1788) );
  nor2_1 U1981 ( .ip1(n1788), .ip2(n2108), .op(n1791) );
  and2_1 U1982 ( .ip1(n1789), .ip2(n2117), .op(n1790) );
  not_ab_or_c_or_d U1983 ( .ip1(n2119), .ip2(n1792), .ip3(n1791), .ip4(n1790), 
        .op(n1799) );
  nor2_1 U1984 ( .ip1(in2[3]), .ip2(n1793), .op(n1794) );
  ab_or_c_or_d U1985 ( .ip1(in2[3]), .ip2(n1962), .ip3(n1794), .ip4(n2100), 
        .op(n1797) );
  nand2_1 U1986 ( .ip1(n2115), .ip2(n1795), .op(n1796) );
  nand4_1 U1987 ( .ip1(n1799), .ip2(n1798), .ip3(n1797), .ip4(n1796), .op(
        n1804) );
  fulladder U1988 ( .a(n1801), .b(in1[0]), .ci(n1800), .co(n1530), .s(n1802)
         );
  nand2_1 U1989 ( .ip1(n1802), .ip2(n2131), .op(n1803) );
  nand3_1 U1990 ( .ip1(n1805), .ip2(n1804), .ip3(n1803), .op(out[0]) );
  inv_1 U1991 ( .ip(n1806), .op(n1838) );
  nand2_1 U1992 ( .ip1(n2048), .ip2(n1830), .op(n1809) );
  nand2_1 U1993 ( .ip1(n2106), .ip2(n1807), .op(n1808) );
  nand4_1 U1994 ( .ip1(n1811), .ip2(n1810), .ip3(n1809), .ip4(n1808), .op(
        n1812) );
  nand2_1 U1995 ( .ip1(n2014), .ip2(n1812), .op(n1818) );
  nand2_1 U1996 ( .ip1(n1813), .ip2(n1946), .op(n1817) );
  or2_1 U1997 ( .ip1(n1815), .ip2(n1814), .op(n1816) );
  nand3_1 U1998 ( .ip1(n1818), .ip2(n1817), .ip3(n1816), .op(n1819) );
  not_ab_or_c_or_d U1999 ( .ip1(n1820), .ip2(n2022), .ip3(n1854), .ip4(n1819), 
        .op(n1837) );
  nor2_1 U2000 ( .ip1(n1822), .ip2(n1821), .op(n1824) );
  nor3_1 U2001 ( .ip1(n1131), .ip2(n1989), .ip3(n1830), .op(n1823) );
  not_ab_or_c_or_d U2002 ( .ip1(n2096), .ip2(n1825), .ip3(n1824), .ip4(n1823), 
        .op(n1835) );
  fulladder U2003 ( .a(in1[3]), .b(n1827), .ci(n1826), .co(n1455), .s(n1828)
         );
  nand2_1 U2004 ( .ip1(n1828), .ip2(n2131), .op(n1834) );
  nand2_1 U2005 ( .ip1(n1874), .ip2(n1829), .op(n1833) );
  nand2_1 U2006 ( .ip1(n1131), .ip2(n1830), .op(n1831) );
  nand2_1 U2007 ( .ip1(n2099), .ip2(n1831), .op(n1832) );
  nand4_1 U2008 ( .ip1(n1835), .ip2(n1834), .ip3(n1833), .ip4(n1832), .op(
        n1836) );
  ab_or_c_or_d U2009 ( .ip1(n1839), .ip2(n1838), .ip3(n1837), .ip4(n1836), 
        .op(out[3]) );
  nor2_1 U2010 ( .ip1(n1841), .ip2(n1840), .op(n1872) );
  nor2_1 U2011 ( .ip1(n1843), .ip2(n1842), .op(n1844) );
  nor2_1 U2012 ( .ip1(n1845), .ip2(n1844), .op(n1846) );
  nor2_1 U2013 ( .ip1(n1847), .ip2(n1846), .op(n1871) );
  nor2_1 U2014 ( .ip1(n1941), .ip2(n1848), .op(n1851) );
  nor2_1 U2015 ( .ip1(n2003), .ip2(n1849), .op(n1850) );
  ab_or_c_or_d U2016 ( .ip1(n1852), .ip2(n2015), .ip3(n1851), .ip4(n1850), 
        .op(n1853) );
  not_ab_or_c_or_d U2017 ( .ip1(n1855), .ip2(n2014), .ip3(n1854), .ip4(n1853), 
        .op(n1870) );
  nor2_1 U2018 ( .ip1(in2[5]), .ip2(in1[5]), .op(n1856) );
  nor2_1 U2019 ( .ip1(n1856), .ip2(n2046), .op(n1860) );
  inv_1 U2020 ( .ip(in2[5]), .op(n1858) );
  nor3_1 U2021 ( .ip1(n1989), .ip2(n1858), .ip3(n1857), .op(n1859) );
  not_ab_or_c_or_d U2022 ( .ip1(n2096), .ip2(n1861), .ip3(n1860), .ip4(n1859), 
        .op(n1868) );
  fulladder U2023 ( .a(in1[5]), .b(n1863), .ci(n1862), .co(n1425), .s(n1864)
         );
  nand2_1 U2024 ( .ip1(n1864), .ip2(n2131), .op(n1867) );
  nand2_1 U2025 ( .ip1(n1876), .ip2(n1865), .op(n1866) );
  nand3_1 U2026 ( .ip1(n1868), .ip2(n1867), .ip3(n1866), .op(n1869) );
  or4_1 U2027 ( .ip1(n1872), .ip2(n1871), .ip3(n1870), .ip4(n1869), .op(out[5]) );
  nand2_1 U2028 ( .ip1(n1874), .ip2(n1873), .op(n1878) );
  nand2_1 U2029 ( .ip1(n1876), .ip2(n1875), .op(n1877) );
  nand2_1 U2030 ( .ip1(n1878), .ip2(n1877), .op(n1903) );
  nor2_1 U2031 ( .ip1(n1985), .ip2(in1[14]), .op(n1879) );
  not_ab_or_c_or_d U2032 ( .ip1(n2092), .ip2(in1[14]), .ip3(n1879), .ip4(n2099), .op(n1881) );
  nor2_1 U2033 ( .ip1(n1881), .ip2(n1880), .op(n1884) );
  nor2_1 U2034 ( .ip1(n2046), .ip2(n1882), .op(n1883) );
  not_ab_or_c_or_d U2035 ( .ip1(n2096), .ip2(n1885), .ip3(n1884), .ip4(n1883), 
        .op(n1900) );
  or2_1 U2036 ( .ip1(n1886), .ip2(n1907), .op(n1899) );
  nor2_1 U2037 ( .ip1(n1131), .ip2(n1887), .op(n1890) );
  nor2_1 U2038 ( .ip1(n1941), .ip2(n1888), .op(n1889) );
  not_ab_or_c_or_d U2039 ( .ip1(n1891), .ip2(n2014), .ip3(n1890), .ip4(n1889), 
        .op(n1892) );
  nand2_1 U2040 ( .ip1(n1893), .ip2(n1892), .op(n1898) );
  fulladder U2041 ( .a(in1[14]), .b(n1895), .ci(n1894), .co(n1184), .s(n1896)
         );
  nand2_1 U2042 ( .ip1(n1896), .ip2(n2131), .op(n1897) );
  nand4_1 U2043 ( .ip1(n1900), .ip2(n1899), .ip3(n1898), .ip4(n1897), .op(
        n1901) );
  ab_or_c_or_d U2044 ( .ip1(n2014), .ip2(n1903), .ip3(n1902), .ip4(n1901), 
        .op(out[14]) );
  nor2_1 U2045 ( .ip1(n1904), .ip2(n1149), .op(n1905) );
  not_ab_or_c_or_d U2046 ( .ip1(n1906), .ip2(n1149), .ip3(n1131), .ip4(n1905), 
        .op(n1908) );
  not_ab_or_c_or_d U2047 ( .ip1(n1909), .ip2(n1131), .ip3(n1908), .ip4(n1907), 
        .op(n1921) );
  nor2_1 U2048 ( .ip1(in2[18]), .ip2(in1[18]), .op(n1910) );
  nor2_1 U2049 ( .ip1(n1910), .ip2(n2046), .op(n1919) );
  nor2_1 U2050 ( .ip1(n1911), .ip2(n1985), .op(n1918) );
  nor2_1 U2051 ( .ip1(n1913), .ip2(n1912), .op(n1917) );
  nor3_1 U2052 ( .ip1(n1989), .ip2(n1915), .ip3(n1914), .op(n1916) );
  or4_1 U2053 ( .ip1(n1919), .ip2(n1918), .ip3(n1917), .ip4(n1916), .op(n1920)
         );
  not_ab_or_c_or_d U2054 ( .ip1(n1923), .ip2(n1922), .ip3(n1921), .ip4(n1920), 
        .op(n1932) );
  fulladder U2055 ( .a(in1[18]), .b(n1925), .ci(n1924), .co(n1096), .s(n1930)
         );
  nor2_1 U2056 ( .ip1(n1927), .ip2(n1926), .op(n1929) );
  not_ab_or_c_or_d U2057 ( .ip1(n1930), .ip2(n2131), .ip3(n1929), .ip4(n1928), 
        .op(n1931) );
  nand2_1 U2058 ( .ip1(n1932), .ip2(n1931), .op(out[18]) );
  fulladder U2059 ( .a(in1[24]), .b(n1934), .ci(n1933), .co(n926), .s(n1959)
         );
  nand2_1 U2060 ( .ip1(n1936), .ip2(n1935), .op(n1940) );
  nand2_1 U2061 ( .ip1(n1938), .ip2(n1937), .op(n1939) );
  nand2_1 U2062 ( .ip1(n1940), .ip2(n1939), .op(n2021) );
  nor2_1 U2063 ( .ip1(n2024), .ip2(n2021), .op(n1944) );
  nor2_1 U2064 ( .ip1(n1941), .ip2(n2016), .op(n1942) );
  ab_or_c_or_d U2065 ( .ip1(n2015), .ip2(n2004), .ip3(in2[4]), .ip4(n1942), 
        .op(n1943) );
  not_ab_or_c_or_d U2066 ( .ip1(n1946), .ip2(n1945), .ip3(n1944), .ip4(n1943), 
        .op(n1950) );
  nor2_1 U2067 ( .ip1(n1947), .ip2(n1978), .op(n1948) );
  nor2_1 U2068 ( .ip1(n2037), .ip2(n1948), .op(n1949) );
  nor2_1 U2069 ( .ip1(n1950), .ip2(n1949), .op(n1958) );
  or2_1 U2070 ( .ip1(in2[24]), .ip2(in1[24]), .op(n1956) );
  nor2_1 U2071 ( .ip1(n1951), .ip2(n1985), .op(n1955) );
  inv_1 U2072 ( .ip(in2[24]), .op(n1953) );
  nor3_1 U2073 ( .ip1(n1989), .ip2(n1953), .ip3(n1952), .op(n1954) );
  ab_or_c_or_d U2074 ( .ip1(n2099), .ip2(n1956), .ip3(n1955), .ip4(n1954), 
        .op(n1957) );
  not_ab_or_c_or_d U2075 ( .ip1(n1959), .ip2(n2131), .ip3(n1958), .ip4(n1957), 
        .op(n1965) );
  nand2_1 U2076 ( .ip1(n1960), .ip2(n2027), .op(n1961) );
  nand2_1 U2077 ( .ip1(n1962), .ip2(n1961), .op(n1963) );
  nand3_1 U2078 ( .ip1(n1965), .ip2(n1964), .ip3(n1963), .op(out[24]) );
  fulladder U2079 ( .a(in1[27]), .b(n1967), .ci(n1966), .co(n2038), .s(n1996)
         );
  inv_1 U2080 ( .ip(n2115), .op(n2053) );
  nor2_1 U2081 ( .ip1(n2053), .ip2(n2116), .op(n1977) );
  nand4_1 U2082 ( .ip1(n1971), .ip2(n1970), .ip3(n1969), .ip4(n1968), .op(
        n2114) );
  nor2_1 U2083 ( .ip1(n2108), .ip2(n2114), .op(n1976) );
  inv_1 U2084 ( .ip(n2119), .op(n1973) );
  nor2_1 U2085 ( .ip1(n1973), .ip2(n1972), .op(n1975) );
  inv_1 U2086 ( .ip(n2117), .op(n2061) );
  nor2_1 U2087 ( .ip1(n2061), .ip2(n2118), .op(n1974) );
  or4_1 U2088 ( .ip1(n1977), .ip2(n1976), .ip3(n1975), .ip4(n1974), .op(n1982)
         );
  nor2_1 U2089 ( .ip1(n1979), .ip2(n1978), .op(n1980) );
  nor2_1 U2090 ( .ip1(n2037), .ip2(n1980), .op(n1981) );
  nor2_1 U2091 ( .ip1(n1982), .ip2(n1981), .op(n1995) );
  nor2_1 U2092 ( .ip1(n1983), .ip2(n2027), .op(n1993) );
  nor2_1 U2093 ( .ip1(in2[27]), .ip2(in1[27]), .op(n1984) );
  nor2_1 U2094 ( .ip1(n1984), .ip2(n2046), .op(n1992) );
  nor2_1 U2095 ( .ip1(n1986), .ip2(n1985), .op(n1991) );
  nor3_1 U2096 ( .ip1(n1989), .ip2(n1988), .ip3(n1987), .op(n1990) );
  or4_1 U2097 ( .ip1(n1993), .ip2(n1992), .ip3(n1991), .ip4(n1990), .op(n1994)
         );
  not_ab_or_c_or_d U2098 ( .ip1(n1996), .ip2(n2131), .ip3(n1995), .ip4(n1994), 
        .op(n2002) );
  or2_1 U2099 ( .ip1(n2075), .ip2(n1997), .op(n1998) );
  nand2_1 U2100 ( .ip1(n1999), .ip2(n1998), .op(n2000) );
  nand3_1 U2101 ( .ip1(n2002), .ip2(n2001), .ip3(n2000), .op(out[27]) );
  nor2_1 U2102 ( .ip1(n2004), .ip2(n2003), .op(n2020) );
  nand2_1 U2103 ( .ip1(n2006), .ip2(n2005), .op(n2012) );
  or2_1 U2104 ( .ip1(in1[28]), .ip2(in2[1]), .op(n2008) );
  nand2_1 U2105 ( .ip1(n2008), .ip2(n2007), .op(n2010) );
  nand2_1 U2106 ( .ip1(n2010), .ip2(n2009), .op(n2011) );
  nand2_1 U2107 ( .ip1(n2012), .ip2(n2011), .op(n2013) );
  nand2_1 U2108 ( .ip1(n2014), .ip2(n2013), .op(n2018) );
  nand2_1 U2109 ( .ip1(n2016), .ip2(n2015), .op(n2017) );
  nand2_1 U2110 ( .ip1(n2018), .ip2(n2017), .op(n2019) );
  not_ab_or_c_or_d U2111 ( .ip1(n2022), .ip2(n2021), .ip3(n2020), .ip4(n2019), 
        .op(n2036) );
  not_ab_or_c_or_d U2112 ( .ip1(N316), .ip2(n2024), .ip3(in2[4]), .ip4(n2023), 
        .op(n2025) );
  nor2_1 U2113 ( .ip1(n2025), .ip2(n2077), .op(n2035) );
  nand2_1 U2114 ( .ip1(n2096), .ip2(n2026), .op(n2033) );
  nand3_1 U2115 ( .ip1(n2092), .ip2(in1[28]), .ip3(in2[28]), .op(n2032) );
  inv_1 U2116 ( .ip(n2027), .op(n2074) );
  nand2_1 U2117 ( .ip1(n2028), .ip2(n2074), .op(n2031) );
  or2_1 U2118 ( .ip1(in1[28]), .ip2(in2[28]), .op(n2029) );
  nand2_1 U2119 ( .ip1(n2099), .ip2(n2029), .op(n2030) );
  nand4_1 U2120 ( .ip1(n2033), .ip2(n2032), .ip3(n2031), .ip4(n2030), .op(
        n2034) );
  not_ab_or_c_or_d U2121 ( .ip1(n2037), .ip2(n2036), .ip3(n2035), .ip4(n2034), 
        .op(n2045) );
  fulladder U2122 ( .a(in1[28]), .b(n2039), .ci(n2038), .co(n2079), .s(n2040)
         );
  nand2_1 U2123 ( .ip1(n2040), .ip2(n2131), .op(n2044) );
  or2_1 U2124 ( .ip1(n2042), .ip2(n2041), .op(n2043) );
  nand3_1 U2125 ( .ip1(n2045), .ip2(n2044), .ip3(n2043), .op(out[28]) );
  nor2_1 U2126 ( .ip1(in1[29]), .ip2(in2[29]), .op(n2047) );
  nor2_1 U2127 ( .ip1(n2047), .ip2(n2046), .op(n2072) );
  nand2_1 U2128 ( .ip1(in1[29]), .ip2(n2048), .op(n2051) );
  nand4_1 U2129 ( .ip1(n2052), .ip2(n2051), .ip3(n2050), .ip4(n2049), .op(
        n2058) );
  nor2_1 U2130 ( .ip1(n2054), .ip2(n2053), .op(n2057) );
  nor2_1 U2131 ( .ip1(n2055), .ip2(n2100), .op(n2056) );
  not_ab_or_c_or_d U2132 ( .ip1(n2059), .ip2(n2058), .ip3(n2057), .ip4(n2056), 
        .op(n2065) );
  or2_1 U2133 ( .ip1(n2061), .ip2(n2060), .op(n2064) );
  nand2_1 U2134 ( .ip1(n2119), .ip2(n2062), .op(n2063) );
  nand3_1 U2135 ( .ip1(n2065), .ip2(n2064), .ip3(n2063), .op(n2066) );
  nand2_1 U2136 ( .ip1(n2124), .ip2(n2066), .op(n2070) );
  nand2_1 U2137 ( .ip1(n2096), .ip2(n2067), .op(n2069) );
  nand3_1 U2138 ( .ip1(n2092), .ip2(in2[29]), .ip3(in1[29]), .op(n2068) );
  nand3_1 U2139 ( .ip1(n2070), .ip2(n2069), .ip3(n2068), .op(n2071) );
  not_ab_or_c_or_d U2140 ( .ip1(n2074), .ip2(n2073), .ip3(n2072), .ip4(n2071), 
        .op(n2084) );
  not_ab_or_c_or_d U2141 ( .ip1(n2076), .ip2(n1131), .ip3(in2[4]), .ip4(n2075), 
        .op(n2078) );
  or2_1 U2142 ( .ip1(n2078), .ip2(n2077), .op(n2083) );
  fulladder U2143 ( .a(in1[29]), .b(n2080), .ci(n2079), .co(n2087), .s(n2081)
         );
  nand2_1 U2144 ( .ip1(n2081), .ip2(n2131), .op(n2082) );
  nand3_1 U2145 ( .ip1(n2084), .ip2(n2083), .ip3(n2082), .op(out[29]) );
  xor2_1 U2146 ( .ip1(n2085), .ip2(in2[31]), .op(n2086) );
  xor2_1 U2147 ( .ip1(n2086), .ip2(N316), .op(n2090) );
  fulladder U2148 ( .a(in1[30]), .b(n2088), .ci(n2087), .co(n2089), .s(n828)
         );
  xor2_1 U2149 ( .ip1(n2090), .ip2(n2089), .op(n2132) );
  not_ab_or_c_or_d U2150 ( .ip1(n2092), .ip2(in2[31]), .ip3(n2091), .ip4(n2099), .op(n2094) );
  nor2_1 U2151 ( .ip1(n2094), .ip2(n2093), .op(n2130) );
  nand2_1 U2152 ( .ip1(n2096), .ip2(n2095), .op(n2128) );
  nand2_1 U2153 ( .ip1(n2098), .ip2(n2097), .op(n2127) );
  nand2_1 U2154 ( .ip1(n2099), .ip2(in2[31]), .op(n2126) );
  nor2_1 U2155 ( .ip1(n2101), .ip2(n2100), .op(n2113) );
  nor2_1 U2156 ( .ip1(n2103), .ip2(n2102), .op(n2104) );
  not_ab_or_c_or_d U2157 ( .ip1(n2106), .ip2(in1[30]), .ip3(n2105), .ip4(n2104), .op(n2107) );
  or2_1 U2158 ( .ip1(n2107), .ip2(n2108), .op(n2111) );
  or2_1 U2159 ( .ip1(n2109), .ip2(n2108), .op(n2110) );
  nand2_1 U2160 ( .ip1(n2111), .ip2(n2110), .op(n2112) );
  not_ab_or_c_or_d U2161 ( .ip1(n2115), .ip2(n2114), .ip3(n2113), .ip4(n2112), 
        .op(n2122) );
  nand2_1 U2162 ( .ip1(n2117), .ip2(n2116), .op(n2121) );
  nand2_1 U2163 ( .ip1(n2119), .ip2(n2118), .op(n2120) );
  nand3_1 U2164 ( .ip1(n2122), .ip2(n2121), .ip3(n2120), .op(n2123) );
  nand2_1 U2165 ( .ip1(n2124), .ip2(n2123), .op(n2125) );
  nand4_1 U2166 ( .ip1(n2128), .ip2(n2127), .ip3(n2126), .ip4(n2125), .op(
        n2129) );
  ab_or_c_or_d U2167 ( .ip1(n2132), .ip2(n2131), .ip3(n2130), .ip4(n2129), 
        .op(out[31]) );
endmodule

