
module vscale_core ( clk, ext_interrupts, imem_haddr, imem_hwrite, imem_hsize, 
        imem_hburst, imem_hmastlock, imem_hprot, imem_htrans, imem_hwdata, 
        imem_hrdata, imem_hready, imem_hresp, dmem_haddr, dmem_hwrite, 
        dmem_hsize, dmem_hburst, dmem_hmastlock, dmem_hprot, dmem_htrans, 
        dmem_hwdata, dmem_hrdata, dmem_hready, dmem_hresp, htif_reset, htif_id, 
        htif_pcr_req_valid, htif_pcr_req_ready, htif_pcr_req_rw, 
        htif_pcr_req_addr, htif_pcr_req_data, htif_pcr_resp_valid, 
        htif_pcr_resp_ready, htif_pcr_resp_data, htif_ipi_req_ready, 
        htif_ipi_req_valid, htif_ipi_req_data, htif_ipi_resp_ready, 
        htif_ipi_resp_valid, htif_ipi_resp_data, htif_debug_stats_pcr );
  input [23:0] ext_interrupts;
  output [31:0] imem_haddr;
  output [2:0] imem_hsize;
  output [2:0] imem_hburst;
  output [3:0] imem_hprot;
  output [1:0] imem_htrans;
  output [31:0] imem_hwdata;
  input [31:0] imem_hrdata;
  input [0:0] imem_hresp;
  output [31:0] dmem_haddr;
  output [2:0] dmem_hsize;
  output [2:0] dmem_hburst;
  output [3:0] dmem_hprot;
  output [1:0] dmem_htrans;
  output [31:0] dmem_hwdata;
  input [31:0] dmem_hrdata;
  input [0:0] dmem_hresp;
  input [11:0] htif_pcr_req_addr;
  input [63:0] htif_pcr_req_data;
  output [63:0] htif_pcr_resp_data;
  input clk, imem_hready, dmem_hready, htif_reset, htif_id, htif_pcr_req_valid,
         htif_pcr_req_rw, htif_pcr_resp_ready, htif_ipi_req_ready,
         htif_ipi_resp_valid, htif_ipi_resp_data;
  output imem_hwrite, imem_hmastlock, dmem_hwrite, dmem_hmastlock,
         htif_pcr_req_ready, htif_pcr_resp_valid, htif_ipi_req_valid,
         htif_ipi_req_data, htif_ipi_resp_ready, htif_debug_stats_pcr;
  wire   imem_badmem_e, dmem_badmem_e, \pipeline/imm[31] ,
         \pipeline/dmem_type[2] , \pipeline/ctrl/wfi_unkilled_WB ,
         \pipeline/ctrl/uses_md_WB , \pipeline/ctrl/dmem_en_WB ,
         \pipeline/ctrl/wr_reg_unkilled_WB , \pipeline/ctrl/had_ex_WB ,
         \pipeline/ctrl/prev_killed_WB , \pipeline/ctrl/prev_killed_DX ,
         \pipeline/ctrl/had_ex_DX , \pipeline/ctrl/N66 ,
         \pipeline/ctrl/store_in_WB , \pipeline/ctrl/replay_IF ,
         \pipeline/regfile/data[31][31] , \pipeline/regfile/data[31][30] ,
         \pipeline/regfile/data[31][29] , \pipeline/regfile/data[31][28] ,
         \pipeline/regfile/data[31][27] , \pipeline/regfile/data[31][26] ,
         \pipeline/regfile/data[31][25] , \pipeline/regfile/data[31][24] ,
         \pipeline/regfile/data[31][23] , \pipeline/regfile/data[31][22] ,
         \pipeline/regfile/data[31][21] , \pipeline/regfile/data[31][20] ,
         \pipeline/regfile/data[31][19] , \pipeline/regfile/data[31][18] ,
         \pipeline/regfile/data[31][17] , \pipeline/regfile/data[31][16] ,
         \pipeline/regfile/data[31][15] , \pipeline/regfile/data[31][14] ,
         \pipeline/regfile/data[31][13] , \pipeline/regfile/data[31][12] ,
         \pipeline/regfile/data[31][11] , \pipeline/regfile/data[31][10] ,
         \pipeline/regfile/data[31][9] , \pipeline/regfile/data[31][8] ,
         \pipeline/regfile/data[31][7] , \pipeline/regfile/data[31][6] ,
         \pipeline/regfile/data[31][5] , \pipeline/regfile/data[31][4] ,
         \pipeline/regfile/data[31][3] , \pipeline/regfile/data[31][2] ,
         \pipeline/regfile/data[31][1] , \pipeline/regfile/data[31][0] ,
         \pipeline/regfile/data[30][31] , \pipeline/regfile/data[30][30] ,
         \pipeline/regfile/data[30][29] , \pipeline/regfile/data[30][28] ,
         \pipeline/regfile/data[30][27] , \pipeline/regfile/data[30][26] ,
         \pipeline/regfile/data[30][25] , \pipeline/regfile/data[30][24] ,
         \pipeline/regfile/data[30][23] , \pipeline/regfile/data[30][22] ,
         \pipeline/regfile/data[30][21] , \pipeline/regfile/data[30][20] ,
         \pipeline/regfile/data[30][19] , \pipeline/regfile/data[30][18] ,
         \pipeline/regfile/data[30][17] , \pipeline/regfile/data[30][16] ,
         \pipeline/regfile/data[30][15] , \pipeline/regfile/data[30][14] ,
         \pipeline/regfile/data[30][13] , \pipeline/regfile/data[30][12] ,
         \pipeline/regfile/data[30][11] , \pipeline/regfile/data[30][10] ,
         \pipeline/regfile/data[30][9] , \pipeline/regfile/data[30][8] ,
         \pipeline/regfile/data[30][7] , \pipeline/regfile/data[30][6] ,
         \pipeline/regfile/data[30][5] , \pipeline/regfile/data[30][4] ,
         \pipeline/regfile/data[30][3] , \pipeline/regfile/data[30][2] ,
         \pipeline/regfile/data[30][1] , \pipeline/regfile/data[30][0] ,
         \pipeline/regfile/data[29][31] , \pipeline/regfile/data[29][30] ,
         \pipeline/regfile/data[29][29] , \pipeline/regfile/data[29][28] ,
         \pipeline/regfile/data[29][27] , \pipeline/regfile/data[29][26] ,
         \pipeline/regfile/data[29][25] , \pipeline/regfile/data[29][24] ,
         \pipeline/regfile/data[29][23] , \pipeline/regfile/data[29][22] ,
         \pipeline/regfile/data[29][21] , \pipeline/regfile/data[29][20] ,
         \pipeline/regfile/data[29][19] , \pipeline/regfile/data[29][18] ,
         \pipeline/regfile/data[29][17] , \pipeline/regfile/data[29][16] ,
         \pipeline/regfile/data[29][15] , \pipeline/regfile/data[29][14] ,
         \pipeline/regfile/data[29][13] , \pipeline/regfile/data[29][12] ,
         \pipeline/regfile/data[29][11] , \pipeline/regfile/data[29][10] ,
         \pipeline/regfile/data[29][9] , \pipeline/regfile/data[29][8] ,
         \pipeline/regfile/data[29][7] , \pipeline/regfile/data[29][6] ,
         \pipeline/regfile/data[29][5] , \pipeline/regfile/data[29][4] ,
         \pipeline/regfile/data[29][3] , \pipeline/regfile/data[29][2] ,
         \pipeline/regfile/data[29][1] , \pipeline/regfile/data[29][0] ,
         \pipeline/regfile/data[28][31] , \pipeline/regfile/data[28][30] ,
         \pipeline/regfile/data[28][29] , \pipeline/regfile/data[28][28] ,
         \pipeline/regfile/data[28][27] , \pipeline/regfile/data[28][26] ,
         \pipeline/regfile/data[28][25] , \pipeline/regfile/data[28][24] ,
         \pipeline/regfile/data[28][23] , \pipeline/regfile/data[28][22] ,
         \pipeline/regfile/data[28][21] , \pipeline/regfile/data[28][20] ,
         \pipeline/regfile/data[28][19] , \pipeline/regfile/data[28][18] ,
         \pipeline/regfile/data[28][17] , \pipeline/regfile/data[28][16] ,
         \pipeline/regfile/data[28][15] , \pipeline/regfile/data[28][14] ,
         \pipeline/regfile/data[28][13] , \pipeline/regfile/data[28][12] ,
         \pipeline/regfile/data[28][11] , \pipeline/regfile/data[28][10] ,
         \pipeline/regfile/data[28][9] , \pipeline/regfile/data[28][8] ,
         \pipeline/regfile/data[28][7] , \pipeline/regfile/data[28][6] ,
         \pipeline/regfile/data[28][5] , \pipeline/regfile/data[28][4] ,
         \pipeline/regfile/data[28][3] , \pipeline/regfile/data[28][2] ,
         \pipeline/regfile/data[28][1] , \pipeline/regfile/data[28][0] ,
         \pipeline/regfile/data[27][31] , \pipeline/regfile/data[27][30] ,
         \pipeline/regfile/data[27][29] , \pipeline/regfile/data[27][28] ,
         \pipeline/regfile/data[27][27] , \pipeline/regfile/data[27][26] ,
         \pipeline/regfile/data[27][25] , \pipeline/regfile/data[27][24] ,
         \pipeline/regfile/data[27][23] , \pipeline/regfile/data[27][22] ,
         \pipeline/regfile/data[27][21] , \pipeline/regfile/data[27][20] ,
         \pipeline/regfile/data[27][19] , \pipeline/regfile/data[27][18] ,
         \pipeline/regfile/data[27][17] , \pipeline/regfile/data[27][16] ,
         \pipeline/regfile/data[27][15] , \pipeline/regfile/data[27][14] ,
         \pipeline/regfile/data[27][13] , \pipeline/regfile/data[27][12] ,
         \pipeline/regfile/data[27][11] , \pipeline/regfile/data[27][10] ,
         \pipeline/regfile/data[27][9] , \pipeline/regfile/data[27][8] ,
         \pipeline/regfile/data[27][7] , \pipeline/regfile/data[27][6] ,
         \pipeline/regfile/data[27][5] , \pipeline/regfile/data[27][4] ,
         \pipeline/regfile/data[27][3] , \pipeline/regfile/data[27][2] ,
         \pipeline/regfile/data[27][1] , \pipeline/regfile/data[27][0] ,
         \pipeline/regfile/data[26][31] , \pipeline/regfile/data[26][30] ,
         \pipeline/regfile/data[26][29] , \pipeline/regfile/data[26][28] ,
         \pipeline/regfile/data[26][27] , \pipeline/regfile/data[26][26] ,
         \pipeline/regfile/data[26][25] , \pipeline/regfile/data[26][24] ,
         \pipeline/regfile/data[26][23] , \pipeline/regfile/data[26][22] ,
         \pipeline/regfile/data[26][21] , \pipeline/regfile/data[26][20] ,
         \pipeline/regfile/data[26][19] , \pipeline/regfile/data[26][18] ,
         \pipeline/regfile/data[26][17] , \pipeline/regfile/data[26][16] ,
         \pipeline/regfile/data[26][15] , \pipeline/regfile/data[26][14] ,
         \pipeline/regfile/data[26][13] , \pipeline/regfile/data[26][12] ,
         \pipeline/regfile/data[26][11] , \pipeline/regfile/data[26][10] ,
         \pipeline/regfile/data[26][9] , \pipeline/regfile/data[26][8] ,
         \pipeline/regfile/data[26][7] , \pipeline/regfile/data[26][6] ,
         \pipeline/regfile/data[26][5] , \pipeline/regfile/data[26][4] ,
         \pipeline/regfile/data[26][3] , \pipeline/regfile/data[26][2] ,
         \pipeline/regfile/data[26][1] , \pipeline/regfile/data[26][0] ,
         \pipeline/regfile/data[25][31] , \pipeline/regfile/data[25][30] ,
         \pipeline/regfile/data[25][29] , \pipeline/regfile/data[25][28] ,
         \pipeline/regfile/data[25][27] , \pipeline/regfile/data[25][26] ,
         \pipeline/regfile/data[25][25] , \pipeline/regfile/data[25][24] ,
         \pipeline/regfile/data[25][23] , \pipeline/regfile/data[25][22] ,
         \pipeline/regfile/data[25][21] , \pipeline/regfile/data[25][20] ,
         \pipeline/regfile/data[25][19] , \pipeline/regfile/data[25][18] ,
         \pipeline/regfile/data[25][17] , \pipeline/regfile/data[25][16] ,
         \pipeline/regfile/data[25][15] , \pipeline/regfile/data[25][14] ,
         \pipeline/regfile/data[25][13] , \pipeline/regfile/data[25][12] ,
         \pipeline/regfile/data[25][11] , \pipeline/regfile/data[25][10] ,
         \pipeline/regfile/data[25][9] , \pipeline/regfile/data[25][8] ,
         \pipeline/regfile/data[25][7] , \pipeline/regfile/data[25][6] ,
         \pipeline/regfile/data[25][5] , \pipeline/regfile/data[25][4] ,
         \pipeline/regfile/data[25][3] , \pipeline/regfile/data[25][2] ,
         \pipeline/regfile/data[25][1] , \pipeline/regfile/data[25][0] ,
         \pipeline/regfile/data[24][31] , \pipeline/regfile/data[24][30] ,
         \pipeline/regfile/data[24][29] , \pipeline/regfile/data[24][28] ,
         \pipeline/regfile/data[24][27] , \pipeline/regfile/data[24][26] ,
         \pipeline/regfile/data[24][25] , \pipeline/regfile/data[24][24] ,
         \pipeline/regfile/data[24][23] , \pipeline/regfile/data[24][22] ,
         \pipeline/regfile/data[24][21] , \pipeline/regfile/data[24][20] ,
         \pipeline/regfile/data[24][19] , \pipeline/regfile/data[24][18] ,
         \pipeline/regfile/data[24][17] , \pipeline/regfile/data[24][16] ,
         \pipeline/regfile/data[24][15] , \pipeline/regfile/data[24][14] ,
         \pipeline/regfile/data[24][13] , \pipeline/regfile/data[24][12] ,
         \pipeline/regfile/data[24][11] , \pipeline/regfile/data[24][10] ,
         \pipeline/regfile/data[24][9] , \pipeline/regfile/data[24][8] ,
         \pipeline/regfile/data[24][7] , \pipeline/regfile/data[24][6] ,
         \pipeline/regfile/data[24][5] , \pipeline/regfile/data[24][4] ,
         \pipeline/regfile/data[24][3] , \pipeline/regfile/data[24][2] ,
         \pipeline/regfile/data[24][1] , \pipeline/regfile/data[24][0] ,
         \pipeline/regfile/data[23][31] , \pipeline/regfile/data[23][30] ,
         \pipeline/regfile/data[23][29] , \pipeline/regfile/data[23][28] ,
         \pipeline/regfile/data[23][27] , \pipeline/regfile/data[23][26] ,
         \pipeline/regfile/data[23][25] , \pipeline/regfile/data[23][24] ,
         \pipeline/regfile/data[23][23] , \pipeline/regfile/data[23][22] ,
         \pipeline/regfile/data[23][21] , \pipeline/regfile/data[23][20] ,
         \pipeline/regfile/data[23][19] , \pipeline/regfile/data[23][18] ,
         \pipeline/regfile/data[23][17] , \pipeline/regfile/data[23][16] ,
         \pipeline/regfile/data[23][15] , \pipeline/regfile/data[23][14] ,
         \pipeline/regfile/data[23][13] , \pipeline/regfile/data[23][12] ,
         \pipeline/regfile/data[23][11] , \pipeline/regfile/data[23][10] ,
         \pipeline/regfile/data[23][9] , \pipeline/regfile/data[23][8] ,
         \pipeline/regfile/data[23][7] , \pipeline/regfile/data[23][6] ,
         \pipeline/regfile/data[23][5] , \pipeline/regfile/data[23][4] ,
         \pipeline/regfile/data[23][3] , \pipeline/regfile/data[23][2] ,
         \pipeline/regfile/data[23][1] , \pipeline/regfile/data[23][0] ,
         \pipeline/regfile/data[22][31] , \pipeline/regfile/data[22][30] ,
         \pipeline/regfile/data[22][29] , \pipeline/regfile/data[22][28] ,
         \pipeline/regfile/data[22][27] , \pipeline/regfile/data[22][26] ,
         \pipeline/regfile/data[22][25] , \pipeline/regfile/data[22][24] ,
         \pipeline/regfile/data[22][23] , \pipeline/regfile/data[22][22] ,
         \pipeline/regfile/data[22][21] , \pipeline/regfile/data[22][20] ,
         \pipeline/regfile/data[22][19] , \pipeline/regfile/data[22][18] ,
         \pipeline/regfile/data[22][17] , \pipeline/regfile/data[22][16] ,
         \pipeline/regfile/data[22][15] , \pipeline/regfile/data[22][14] ,
         \pipeline/regfile/data[22][13] , \pipeline/regfile/data[22][12] ,
         \pipeline/regfile/data[22][11] , \pipeline/regfile/data[22][10] ,
         \pipeline/regfile/data[22][9] , \pipeline/regfile/data[22][8] ,
         \pipeline/regfile/data[22][7] , \pipeline/regfile/data[22][6] ,
         \pipeline/regfile/data[22][5] , \pipeline/regfile/data[22][4] ,
         \pipeline/regfile/data[22][3] , \pipeline/regfile/data[22][2] ,
         \pipeline/regfile/data[22][1] , \pipeline/regfile/data[22][0] ,
         \pipeline/regfile/data[21][31] , \pipeline/regfile/data[21][30] ,
         \pipeline/regfile/data[21][29] , \pipeline/regfile/data[21][28] ,
         \pipeline/regfile/data[21][27] , \pipeline/regfile/data[21][26] ,
         \pipeline/regfile/data[21][25] , \pipeline/regfile/data[21][24] ,
         \pipeline/regfile/data[21][23] , \pipeline/regfile/data[21][22] ,
         \pipeline/regfile/data[21][21] , \pipeline/regfile/data[21][20] ,
         \pipeline/regfile/data[21][19] , \pipeline/regfile/data[21][18] ,
         \pipeline/regfile/data[21][17] , \pipeline/regfile/data[21][16] ,
         \pipeline/regfile/data[21][15] , \pipeline/regfile/data[21][14] ,
         \pipeline/regfile/data[21][13] , \pipeline/regfile/data[21][12] ,
         \pipeline/regfile/data[21][11] , \pipeline/regfile/data[21][10] ,
         \pipeline/regfile/data[21][9] , \pipeline/regfile/data[21][8] ,
         \pipeline/regfile/data[21][7] , \pipeline/regfile/data[21][6] ,
         \pipeline/regfile/data[21][5] , \pipeline/regfile/data[21][4] ,
         \pipeline/regfile/data[21][3] , \pipeline/regfile/data[21][2] ,
         \pipeline/regfile/data[21][1] , \pipeline/regfile/data[21][0] ,
         \pipeline/regfile/data[20][31] , \pipeline/regfile/data[20][30] ,
         \pipeline/regfile/data[20][29] , \pipeline/regfile/data[20][28] ,
         \pipeline/regfile/data[20][27] , \pipeline/regfile/data[20][26] ,
         \pipeline/regfile/data[20][25] , \pipeline/regfile/data[20][24] ,
         \pipeline/regfile/data[20][23] , \pipeline/regfile/data[20][22] ,
         \pipeline/regfile/data[20][21] , \pipeline/regfile/data[20][20] ,
         \pipeline/regfile/data[20][19] , \pipeline/regfile/data[20][18] ,
         \pipeline/regfile/data[20][17] , \pipeline/regfile/data[20][16] ,
         \pipeline/regfile/data[20][15] , \pipeline/regfile/data[20][14] ,
         \pipeline/regfile/data[20][13] , \pipeline/regfile/data[20][12] ,
         \pipeline/regfile/data[20][11] , \pipeline/regfile/data[20][10] ,
         \pipeline/regfile/data[20][9] , \pipeline/regfile/data[20][8] ,
         \pipeline/regfile/data[20][7] , \pipeline/regfile/data[20][6] ,
         \pipeline/regfile/data[20][5] , \pipeline/regfile/data[20][4] ,
         \pipeline/regfile/data[20][3] , \pipeline/regfile/data[20][2] ,
         \pipeline/regfile/data[20][1] , \pipeline/regfile/data[20][0] ,
         \pipeline/regfile/data[19][31] , \pipeline/regfile/data[19][30] ,
         \pipeline/regfile/data[19][29] , \pipeline/regfile/data[19][28] ,
         \pipeline/regfile/data[19][27] , \pipeline/regfile/data[19][26] ,
         \pipeline/regfile/data[19][25] , \pipeline/regfile/data[19][24] ,
         \pipeline/regfile/data[19][23] , \pipeline/regfile/data[19][22] ,
         \pipeline/regfile/data[19][21] , \pipeline/regfile/data[19][20] ,
         \pipeline/regfile/data[19][19] , \pipeline/regfile/data[19][18] ,
         \pipeline/regfile/data[19][17] , \pipeline/regfile/data[19][16] ,
         \pipeline/regfile/data[19][15] , \pipeline/regfile/data[19][14] ,
         \pipeline/regfile/data[19][13] , \pipeline/regfile/data[19][12] ,
         \pipeline/regfile/data[19][11] , \pipeline/regfile/data[19][10] ,
         \pipeline/regfile/data[19][9] , \pipeline/regfile/data[19][8] ,
         \pipeline/regfile/data[19][7] , \pipeline/regfile/data[19][6] ,
         \pipeline/regfile/data[19][5] , \pipeline/regfile/data[19][4] ,
         \pipeline/regfile/data[19][3] , \pipeline/regfile/data[19][2] ,
         \pipeline/regfile/data[19][1] , \pipeline/regfile/data[19][0] ,
         \pipeline/regfile/data[18][31] , \pipeline/regfile/data[18][30] ,
         \pipeline/regfile/data[18][29] , \pipeline/regfile/data[18][28] ,
         \pipeline/regfile/data[18][27] , \pipeline/regfile/data[18][26] ,
         \pipeline/regfile/data[18][25] , \pipeline/regfile/data[18][24] ,
         \pipeline/regfile/data[18][23] , \pipeline/regfile/data[18][22] ,
         \pipeline/regfile/data[18][21] , \pipeline/regfile/data[18][20] ,
         \pipeline/regfile/data[18][19] , \pipeline/regfile/data[18][18] ,
         \pipeline/regfile/data[18][17] , \pipeline/regfile/data[18][16] ,
         \pipeline/regfile/data[18][15] , \pipeline/regfile/data[18][14] ,
         \pipeline/regfile/data[18][13] , \pipeline/regfile/data[18][12] ,
         \pipeline/regfile/data[18][11] , \pipeline/regfile/data[18][10] ,
         \pipeline/regfile/data[18][9] , \pipeline/regfile/data[18][8] ,
         \pipeline/regfile/data[18][7] , \pipeline/regfile/data[18][6] ,
         \pipeline/regfile/data[18][5] , \pipeline/regfile/data[18][4] ,
         \pipeline/regfile/data[18][3] , \pipeline/regfile/data[18][2] ,
         \pipeline/regfile/data[18][1] , \pipeline/regfile/data[18][0] ,
         \pipeline/regfile/data[17][31] , \pipeline/regfile/data[17][30] ,
         \pipeline/regfile/data[17][29] , \pipeline/regfile/data[17][28] ,
         \pipeline/regfile/data[17][27] , \pipeline/regfile/data[17][26] ,
         \pipeline/regfile/data[17][25] , \pipeline/regfile/data[17][24] ,
         \pipeline/regfile/data[17][23] , \pipeline/regfile/data[17][22] ,
         \pipeline/regfile/data[17][21] , \pipeline/regfile/data[17][20] ,
         \pipeline/regfile/data[17][19] , \pipeline/regfile/data[17][18] ,
         \pipeline/regfile/data[17][17] , \pipeline/regfile/data[17][16] ,
         \pipeline/regfile/data[17][15] , \pipeline/regfile/data[17][14] ,
         \pipeline/regfile/data[17][13] , \pipeline/regfile/data[17][12] ,
         \pipeline/regfile/data[17][11] , \pipeline/regfile/data[17][10] ,
         \pipeline/regfile/data[17][9] , \pipeline/regfile/data[17][8] ,
         \pipeline/regfile/data[17][7] , \pipeline/regfile/data[17][6] ,
         \pipeline/regfile/data[17][5] , \pipeline/regfile/data[17][4] ,
         \pipeline/regfile/data[17][3] , \pipeline/regfile/data[17][2] ,
         \pipeline/regfile/data[17][1] , \pipeline/regfile/data[17][0] ,
         \pipeline/regfile/data[16][31] , \pipeline/regfile/data[16][30] ,
         \pipeline/regfile/data[16][29] , \pipeline/regfile/data[16][28] ,
         \pipeline/regfile/data[16][27] , \pipeline/regfile/data[16][26] ,
         \pipeline/regfile/data[16][25] , \pipeline/regfile/data[16][24] ,
         \pipeline/regfile/data[16][23] , \pipeline/regfile/data[16][22] ,
         \pipeline/regfile/data[16][21] , \pipeline/regfile/data[16][20] ,
         \pipeline/regfile/data[16][19] , \pipeline/regfile/data[16][18] ,
         \pipeline/regfile/data[16][17] , \pipeline/regfile/data[16][16] ,
         \pipeline/regfile/data[16][15] , \pipeline/regfile/data[16][14] ,
         \pipeline/regfile/data[16][13] , \pipeline/regfile/data[16][12] ,
         \pipeline/regfile/data[16][11] , \pipeline/regfile/data[16][10] ,
         \pipeline/regfile/data[16][9] , \pipeline/regfile/data[16][8] ,
         \pipeline/regfile/data[16][7] , \pipeline/regfile/data[16][6] ,
         \pipeline/regfile/data[16][5] , \pipeline/regfile/data[16][4] ,
         \pipeline/regfile/data[16][3] , \pipeline/regfile/data[16][2] ,
         \pipeline/regfile/data[16][1] , \pipeline/regfile/data[16][0] ,
         \pipeline/regfile/data[15][31] , \pipeline/regfile/data[15][30] ,
         \pipeline/regfile/data[15][29] , \pipeline/regfile/data[15][28] ,
         \pipeline/regfile/data[15][27] , \pipeline/regfile/data[15][26] ,
         \pipeline/regfile/data[15][25] , \pipeline/regfile/data[15][24] ,
         \pipeline/regfile/data[15][23] , \pipeline/regfile/data[15][22] ,
         \pipeline/regfile/data[15][21] , \pipeline/regfile/data[15][20] ,
         \pipeline/regfile/data[15][19] , \pipeline/regfile/data[15][18] ,
         \pipeline/regfile/data[15][17] , \pipeline/regfile/data[15][16] ,
         \pipeline/regfile/data[15][15] , \pipeline/regfile/data[15][14] ,
         \pipeline/regfile/data[15][13] , \pipeline/regfile/data[15][12] ,
         \pipeline/regfile/data[15][11] , \pipeline/regfile/data[15][10] ,
         \pipeline/regfile/data[15][9] , \pipeline/regfile/data[15][8] ,
         \pipeline/regfile/data[15][7] , \pipeline/regfile/data[15][6] ,
         \pipeline/regfile/data[15][5] , \pipeline/regfile/data[15][4] ,
         \pipeline/regfile/data[15][3] , \pipeline/regfile/data[15][2] ,
         \pipeline/regfile/data[15][1] , \pipeline/regfile/data[15][0] ,
         \pipeline/regfile/data[14][31] , \pipeline/regfile/data[14][30] ,
         \pipeline/regfile/data[14][29] , \pipeline/regfile/data[14][28] ,
         \pipeline/regfile/data[14][27] , \pipeline/regfile/data[14][26] ,
         \pipeline/regfile/data[14][25] , \pipeline/regfile/data[14][24] ,
         \pipeline/regfile/data[14][23] , \pipeline/regfile/data[14][22] ,
         \pipeline/regfile/data[14][21] , \pipeline/regfile/data[14][20] ,
         \pipeline/regfile/data[14][19] , \pipeline/regfile/data[14][18] ,
         \pipeline/regfile/data[14][17] , \pipeline/regfile/data[14][16] ,
         \pipeline/regfile/data[14][15] , \pipeline/regfile/data[14][14] ,
         \pipeline/regfile/data[14][13] , \pipeline/regfile/data[14][12] ,
         \pipeline/regfile/data[14][11] , \pipeline/regfile/data[14][10] ,
         \pipeline/regfile/data[14][9] , \pipeline/regfile/data[14][8] ,
         \pipeline/regfile/data[14][7] , \pipeline/regfile/data[14][6] ,
         \pipeline/regfile/data[14][5] , \pipeline/regfile/data[14][4] ,
         \pipeline/regfile/data[14][3] , \pipeline/regfile/data[14][2] ,
         \pipeline/regfile/data[14][1] , \pipeline/regfile/data[14][0] ,
         \pipeline/regfile/data[13][31] , \pipeline/regfile/data[13][30] ,
         \pipeline/regfile/data[13][29] , \pipeline/regfile/data[13][28] ,
         \pipeline/regfile/data[13][27] , \pipeline/regfile/data[13][26] ,
         \pipeline/regfile/data[13][25] , \pipeline/regfile/data[13][24] ,
         \pipeline/regfile/data[13][23] , \pipeline/regfile/data[13][22] ,
         \pipeline/regfile/data[13][21] , \pipeline/regfile/data[13][20] ,
         \pipeline/regfile/data[13][19] , \pipeline/regfile/data[13][18] ,
         \pipeline/regfile/data[13][17] , \pipeline/regfile/data[13][16] ,
         \pipeline/regfile/data[13][15] , \pipeline/regfile/data[13][14] ,
         \pipeline/regfile/data[13][13] , \pipeline/regfile/data[13][12] ,
         \pipeline/regfile/data[13][11] , \pipeline/regfile/data[13][10] ,
         \pipeline/regfile/data[13][9] , \pipeline/regfile/data[13][8] ,
         \pipeline/regfile/data[13][7] , \pipeline/regfile/data[13][6] ,
         \pipeline/regfile/data[13][5] , \pipeline/regfile/data[13][4] ,
         \pipeline/regfile/data[13][3] , \pipeline/regfile/data[13][2] ,
         \pipeline/regfile/data[13][1] , \pipeline/regfile/data[13][0] ,
         \pipeline/regfile/data[12][31] , \pipeline/regfile/data[12][30] ,
         \pipeline/regfile/data[12][29] , \pipeline/regfile/data[12][28] ,
         \pipeline/regfile/data[12][27] , \pipeline/regfile/data[12][26] ,
         \pipeline/regfile/data[12][25] , \pipeline/regfile/data[12][24] ,
         \pipeline/regfile/data[12][23] , \pipeline/regfile/data[12][22] ,
         \pipeline/regfile/data[12][21] , \pipeline/regfile/data[12][20] ,
         \pipeline/regfile/data[12][19] , \pipeline/regfile/data[12][18] ,
         \pipeline/regfile/data[12][17] , \pipeline/regfile/data[12][16] ,
         \pipeline/regfile/data[12][15] , \pipeline/regfile/data[12][14] ,
         \pipeline/regfile/data[12][13] , \pipeline/regfile/data[12][12] ,
         \pipeline/regfile/data[12][11] , \pipeline/regfile/data[12][10] ,
         \pipeline/regfile/data[12][9] , \pipeline/regfile/data[12][8] ,
         \pipeline/regfile/data[12][7] , \pipeline/regfile/data[12][6] ,
         \pipeline/regfile/data[12][5] , \pipeline/regfile/data[12][4] ,
         \pipeline/regfile/data[12][3] , \pipeline/regfile/data[12][2] ,
         \pipeline/regfile/data[12][1] , \pipeline/regfile/data[12][0] ,
         \pipeline/regfile/data[11][31] , \pipeline/regfile/data[11][30] ,
         \pipeline/regfile/data[11][29] , \pipeline/regfile/data[11][28] ,
         \pipeline/regfile/data[11][27] , \pipeline/regfile/data[11][26] ,
         \pipeline/regfile/data[11][25] , \pipeline/regfile/data[11][24] ,
         \pipeline/regfile/data[11][23] , \pipeline/regfile/data[11][22] ,
         \pipeline/regfile/data[11][21] , \pipeline/regfile/data[11][20] ,
         \pipeline/regfile/data[11][19] , \pipeline/regfile/data[11][18] ,
         \pipeline/regfile/data[11][17] , \pipeline/regfile/data[11][16] ,
         \pipeline/regfile/data[11][15] , \pipeline/regfile/data[11][14] ,
         \pipeline/regfile/data[11][13] , \pipeline/regfile/data[11][12] ,
         \pipeline/regfile/data[11][11] , \pipeline/regfile/data[11][10] ,
         \pipeline/regfile/data[11][9] , \pipeline/regfile/data[11][8] ,
         \pipeline/regfile/data[11][7] , \pipeline/regfile/data[11][6] ,
         \pipeline/regfile/data[11][5] , \pipeline/regfile/data[11][4] ,
         \pipeline/regfile/data[11][3] , \pipeline/regfile/data[11][2] ,
         \pipeline/regfile/data[11][1] , \pipeline/regfile/data[11][0] ,
         \pipeline/regfile/data[10][31] , \pipeline/regfile/data[10][30] ,
         \pipeline/regfile/data[10][29] , \pipeline/regfile/data[10][28] ,
         \pipeline/regfile/data[10][27] , \pipeline/regfile/data[10][26] ,
         \pipeline/regfile/data[10][25] , \pipeline/regfile/data[10][24] ,
         \pipeline/regfile/data[10][23] , \pipeline/regfile/data[10][22] ,
         \pipeline/regfile/data[10][21] , \pipeline/regfile/data[10][20] ,
         \pipeline/regfile/data[10][19] , \pipeline/regfile/data[10][18] ,
         \pipeline/regfile/data[10][17] , \pipeline/regfile/data[10][16] ,
         \pipeline/regfile/data[10][15] , \pipeline/regfile/data[10][14] ,
         \pipeline/regfile/data[10][13] , \pipeline/regfile/data[10][12] ,
         \pipeline/regfile/data[10][11] , \pipeline/regfile/data[10][10] ,
         \pipeline/regfile/data[10][9] , \pipeline/regfile/data[10][8] ,
         \pipeline/regfile/data[10][7] , \pipeline/regfile/data[10][6] ,
         \pipeline/regfile/data[10][5] , \pipeline/regfile/data[10][4] ,
         \pipeline/regfile/data[10][3] , \pipeline/regfile/data[10][2] ,
         \pipeline/regfile/data[10][1] , \pipeline/regfile/data[10][0] ,
         \pipeline/regfile/data[9][31] , \pipeline/regfile/data[9][30] ,
         \pipeline/regfile/data[9][29] , \pipeline/regfile/data[9][28] ,
         \pipeline/regfile/data[9][27] , \pipeline/regfile/data[9][26] ,
         \pipeline/regfile/data[9][25] , \pipeline/regfile/data[9][24] ,
         \pipeline/regfile/data[9][23] , \pipeline/regfile/data[9][22] ,
         \pipeline/regfile/data[9][21] , \pipeline/regfile/data[9][20] ,
         \pipeline/regfile/data[9][19] , \pipeline/regfile/data[9][18] ,
         \pipeline/regfile/data[9][17] , \pipeline/regfile/data[9][16] ,
         \pipeline/regfile/data[9][15] , \pipeline/regfile/data[9][14] ,
         \pipeline/regfile/data[9][13] , \pipeline/regfile/data[9][12] ,
         \pipeline/regfile/data[9][11] , \pipeline/regfile/data[9][10] ,
         \pipeline/regfile/data[9][9] , \pipeline/regfile/data[9][8] ,
         \pipeline/regfile/data[9][7] , \pipeline/regfile/data[9][6] ,
         \pipeline/regfile/data[9][5] , \pipeline/regfile/data[9][4] ,
         \pipeline/regfile/data[9][3] , \pipeline/regfile/data[9][2] ,
         \pipeline/regfile/data[9][1] , \pipeline/regfile/data[9][0] ,
         \pipeline/regfile/data[8][31] , \pipeline/regfile/data[8][30] ,
         \pipeline/regfile/data[8][29] , \pipeline/regfile/data[8][28] ,
         \pipeline/regfile/data[8][27] , \pipeline/regfile/data[8][26] ,
         \pipeline/regfile/data[8][25] , \pipeline/regfile/data[8][24] ,
         \pipeline/regfile/data[8][23] , \pipeline/regfile/data[8][22] ,
         \pipeline/regfile/data[8][21] , \pipeline/regfile/data[8][20] ,
         \pipeline/regfile/data[8][19] , \pipeline/regfile/data[8][18] ,
         \pipeline/regfile/data[8][17] , \pipeline/regfile/data[8][16] ,
         \pipeline/regfile/data[8][15] , \pipeline/regfile/data[8][14] ,
         \pipeline/regfile/data[8][13] , \pipeline/regfile/data[8][12] ,
         \pipeline/regfile/data[8][11] , \pipeline/regfile/data[8][10] ,
         \pipeline/regfile/data[8][9] , \pipeline/regfile/data[8][8] ,
         \pipeline/regfile/data[8][7] , \pipeline/regfile/data[8][6] ,
         \pipeline/regfile/data[8][5] , \pipeline/regfile/data[8][4] ,
         \pipeline/regfile/data[8][3] , \pipeline/regfile/data[8][2] ,
         \pipeline/regfile/data[8][1] , \pipeline/regfile/data[8][0] ,
         \pipeline/regfile/data[7][31] , \pipeline/regfile/data[7][30] ,
         \pipeline/regfile/data[7][29] , \pipeline/regfile/data[7][28] ,
         \pipeline/regfile/data[7][27] , \pipeline/regfile/data[7][26] ,
         \pipeline/regfile/data[7][25] , \pipeline/regfile/data[7][24] ,
         \pipeline/regfile/data[7][23] , \pipeline/regfile/data[7][22] ,
         \pipeline/regfile/data[7][21] , \pipeline/regfile/data[7][20] ,
         \pipeline/regfile/data[7][19] , \pipeline/regfile/data[7][18] ,
         \pipeline/regfile/data[7][17] , \pipeline/regfile/data[7][16] ,
         \pipeline/regfile/data[7][15] , \pipeline/regfile/data[7][14] ,
         \pipeline/regfile/data[7][13] , \pipeline/regfile/data[7][12] ,
         \pipeline/regfile/data[7][11] , \pipeline/regfile/data[7][10] ,
         \pipeline/regfile/data[7][9] , \pipeline/regfile/data[7][8] ,
         \pipeline/regfile/data[7][7] , \pipeline/regfile/data[7][6] ,
         \pipeline/regfile/data[7][5] , \pipeline/regfile/data[7][4] ,
         \pipeline/regfile/data[7][3] , \pipeline/regfile/data[7][2] ,
         \pipeline/regfile/data[7][1] , \pipeline/regfile/data[7][0] ,
         \pipeline/regfile/data[6][31] , \pipeline/regfile/data[6][30] ,
         \pipeline/regfile/data[6][29] , \pipeline/regfile/data[6][28] ,
         \pipeline/regfile/data[6][27] , \pipeline/regfile/data[6][26] ,
         \pipeline/regfile/data[6][25] , \pipeline/regfile/data[6][24] ,
         \pipeline/regfile/data[6][23] , \pipeline/regfile/data[6][22] ,
         \pipeline/regfile/data[6][21] , \pipeline/regfile/data[6][20] ,
         \pipeline/regfile/data[6][19] , \pipeline/regfile/data[6][18] ,
         \pipeline/regfile/data[6][17] , \pipeline/regfile/data[6][16] ,
         \pipeline/regfile/data[6][15] , \pipeline/regfile/data[6][14] ,
         \pipeline/regfile/data[6][13] , \pipeline/regfile/data[6][12] ,
         \pipeline/regfile/data[6][11] , \pipeline/regfile/data[6][10] ,
         \pipeline/regfile/data[6][9] , \pipeline/regfile/data[6][8] ,
         \pipeline/regfile/data[6][7] , \pipeline/regfile/data[6][6] ,
         \pipeline/regfile/data[6][5] , \pipeline/regfile/data[6][4] ,
         \pipeline/regfile/data[6][3] , \pipeline/regfile/data[6][2] ,
         \pipeline/regfile/data[6][1] , \pipeline/regfile/data[6][0] ,
         \pipeline/regfile/data[5][31] , \pipeline/regfile/data[5][30] ,
         \pipeline/regfile/data[5][29] , \pipeline/regfile/data[5][28] ,
         \pipeline/regfile/data[5][27] , \pipeline/regfile/data[5][26] ,
         \pipeline/regfile/data[5][25] , \pipeline/regfile/data[5][24] ,
         \pipeline/regfile/data[5][23] , \pipeline/regfile/data[5][22] ,
         \pipeline/regfile/data[5][21] , \pipeline/regfile/data[5][20] ,
         \pipeline/regfile/data[5][19] , \pipeline/regfile/data[5][18] ,
         \pipeline/regfile/data[5][17] , \pipeline/regfile/data[5][16] ,
         \pipeline/regfile/data[5][15] , \pipeline/regfile/data[5][14] ,
         \pipeline/regfile/data[5][13] , \pipeline/regfile/data[5][12] ,
         \pipeline/regfile/data[5][11] , \pipeline/regfile/data[5][10] ,
         \pipeline/regfile/data[5][9] , \pipeline/regfile/data[5][8] ,
         \pipeline/regfile/data[5][7] , \pipeline/regfile/data[5][6] ,
         \pipeline/regfile/data[5][5] , \pipeline/regfile/data[5][4] ,
         \pipeline/regfile/data[5][3] , \pipeline/regfile/data[5][2] ,
         \pipeline/regfile/data[5][1] , \pipeline/regfile/data[5][0] ,
         \pipeline/regfile/data[4][31] , \pipeline/regfile/data[4][30] ,
         \pipeline/regfile/data[4][29] , \pipeline/regfile/data[4][28] ,
         \pipeline/regfile/data[4][27] , \pipeline/regfile/data[4][26] ,
         \pipeline/regfile/data[4][25] , \pipeline/regfile/data[4][24] ,
         \pipeline/regfile/data[4][23] , \pipeline/regfile/data[4][22] ,
         \pipeline/regfile/data[4][21] , \pipeline/regfile/data[4][20] ,
         \pipeline/regfile/data[4][19] , \pipeline/regfile/data[4][18] ,
         \pipeline/regfile/data[4][17] , \pipeline/regfile/data[4][16] ,
         \pipeline/regfile/data[4][15] , \pipeline/regfile/data[4][14] ,
         \pipeline/regfile/data[4][13] , \pipeline/regfile/data[4][12] ,
         \pipeline/regfile/data[4][11] , \pipeline/regfile/data[4][10] ,
         \pipeline/regfile/data[4][9] , \pipeline/regfile/data[4][8] ,
         \pipeline/regfile/data[4][7] , \pipeline/regfile/data[4][6] ,
         \pipeline/regfile/data[4][5] , \pipeline/regfile/data[4][4] ,
         \pipeline/regfile/data[4][3] , \pipeline/regfile/data[4][2] ,
         \pipeline/regfile/data[4][1] , \pipeline/regfile/data[4][0] ,
         \pipeline/regfile/data[3][31] , \pipeline/regfile/data[3][30] ,
         \pipeline/regfile/data[3][29] , \pipeline/regfile/data[3][28] ,
         \pipeline/regfile/data[3][27] , \pipeline/regfile/data[3][26] ,
         \pipeline/regfile/data[3][25] , \pipeline/regfile/data[3][24] ,
         \pipeline/regfile/data[3][23] , \pipeline/regfile/data[3][22] ,
         \pipeline/regfile/data[3][21] , \pipeline/regfile/data[3][20] ,
         \pipeline/regfile/data[3][19] , \pipeline/regfile/data[3][18] ,
         \pipeline/regfile/data[3][17] , \pipeline/regfile/data[3][16] ,
         \pipeline/regfile/data[3][15] , \pipeline/regfile/data[3][14] ,
         \pipeline/regfile/data[3][13] , \pipeline/regfile/data[3][12] ,
         \pipeline/regfile/data[3][11] , \pipeline/regfile/data[3][10] ,
         \pipeline/regfile/data[3][9] , \pipeline/regfile/data[3][8] ,
         \pipeline/regfile/data[3][7] , \pipeline/regfile/data[3][6] ,
         \pipeline/regfile/data[3][5] , \pipeline/regfile/data[3][4] ,
         \pipeline/regfile/data[3][3] , \pipeline/regfile/data[3][2] ,
         \pipeline/regfile/data[3][1] , \pipeline/regfile/data[3][0] ,
         \pipeline/regfile/data[2][31] , \pipeline/regfile/data[2][30] ,
         \pipeline/regfile/data[2][29] , \pipeline/regfile/data[2][28] ,
         \pipeline/regfile/data[2][27] , \pipeline/regfile/data[2][26] ,
         \pipeline/regfile/data[2][25] , \pipeline/regfile/data[2][24] ,
         \pipeline/regfile/data[2][23] , \pipeline/regfile/data[2][22] ,
         \pipeline/regfile/data[2][21] , \pipeline/regfile/data[2][20] ,
         \pipeline/regfile/data[2][19] , \pipeline/regfile/data[2][18] ,
         \pipeline/regfile/data[2][17] , \pipeline/regfile/data[2][16] ,
         \pipeline/regfile/data[2][15] , \pipeline/regfile/data[2][14] ,
         \pipeline/regfile/data[2][13] , \pipeline/regfile/data[2][12] ,
         \pipeline/regfile/data[2][11] , \pipeline/regfile/data[2][10] ,
         \pipeline/regfile/data[2][9] , \pipeline/regfile/data[2][8] ,
         \pipeline/regfile/data[2][7] , \pipeline/regfile/data[2][6] ,
         \pipeline/regfile/data[2][5] , \pipeline/regfile/data[2][4] ,
         \pipeline/regfile/data[2][3] , \pipeline/regfile/data[2][2] ,
         \pipeline/regfile/data[2][1] , \pipeline/regfile/data[2][0] ,
         \pipeline/regfile/data[1][31] , \pipeline/regfile/data[1][30] ,
         \pipeline/regfile/data[1][29] , \pipeline/regfile/data[1][28] ,
         \pipeline/regfile/data[1][27] , \pipeline/regfile/data[1][26] ,
         \pipeline/regfile/data[1][25] , \pipeline/regfile/data[1][24] ,
         \pipeline/regfile/data[1][23] , \pipeline/regfile/data[1][22] ,
         \pipeline/regfile/data[1][21] , \pipeline/regfile/data[1][20] ,
         \pipeline/regfile/data[1][19] , \pipeline/regfile/data[1][18] ,
         \pipeline/regfile/data[1][17] , \pipeline/regfile/data[1][16] ,
         \pipeline/regfile/data[1][15] , \pipeline/regfile/data[1][14] ,
         \pipeline/regfile/data[1][13] , \pipeline/regfile/data[1][12] ,
         \pipeline/regfile/data[1][11] , \pipeline/regfile/data[1][10] ,
         \pipeline/regfile/data[1][9] , \pipeline/regfile/data[1][8] ,
         \pipeline/regfile/data[1][7] , \pipeline/regfile/data[1][6] ,
         \pipeline/regfile/data[1][5] , \pipeline/regfile/data[1][4] ,
         \pipeline/regfile/data[1][3] , \pipeline/regfile/data[1][2] ,
         \pipeline/regfile/data[1][1] , \pipeline/regfile/data[1][0] ,
         \pipeline/md/N162 , \pipeline/md/negate_output , \pipeline/csr/N2387 ,
         \pipeline/csr/N2385 , \pipeline/csr/N2144 , \pipeline/csr/N2143 ,
         \pipeline/csr/N2142 , \pipeline/csr/N2141 , \pipeline/csr/N2140 ,
         \pipeline/csr/N2139 , \pipeline/csr/N2138 , \pipeline/csr/N2137 ,
         \pipeline/csr/N2136 , \pipeline/csr/N2135 , \pipeline/csr/N2134 ,
         \pipeline/csr/N2133 , \pipeline/csr/N2132 , \pipeline/csr/N2131 ,
         \pipeline/csr/N2130 , \pipeline/csr/N2129 , \pipeline/csr/N2128 ,
         \pipeline/csr/N2127 , \pipeline/csr/N2126 , \pipeline/csr/N2125 ,
         \pipeline/csr/N2124 , \pipeline/csr/N2123 , \pipeline/csr/N2122 ,
         \pipeline/csr/N2121 , \pipeline/csr/N2120 , \pipeline/csr/N2119 ,
         \pipeline/csr/N2118 , \pipeline/csr/N2117 , \pipeline/csr/N2116 ,
         \pipeline/csr/N2115 , \pipeline/csr/N2114 , \pipeline/csr/N2113 ,
         \pipeline/csr/N2112 , \pipeline/csr/N2111 , \pipeline/csr/N2110 ,
         \pipeline/csr/N2109 , \pipeline/csr/N2108 , \pipeline/csr/N2107 ,
         \pipeline/csr/N2106 , \pipeline/csr/N2105 , \pipeline/csr/N2104 ,
         \pipeline/csr/N2103 , \pipeline/csr/N2102 , \pipeline/csr/N2101 ,
         \pipeline/csr/N2100 , \pipeline/csr/N2099 , \pipeline/csr/N2098 ,
         \pipeline/csr/N2097 , \pipeline/csr/N2096 , \pipeline/csr/N2095 ,
         \pipeline/csr/N2094 , \pipeline/csr/N2093 , \pipeline/csr/N2092 ,
         \pipeline/csr/N2091 , \pipeline/csr/N2090 , \pipeline/csr/N2089 ,
         \pipeline/csr/N2088 , \pipeline/csr/N2087 , \pipeline/csr/N2086 ,
         \pipeline/csr/N2085 , \pipeline/csr/N2084 , \pipeline/csr/N2083 ,
         \pipeline/csr/N2082 , \pipeline/csr/N2081 , \pipeline/csr/N2000 ,
         \pipeline/csr/N1999 , \pipeline/csr/N1998 , \pipeline/csr/N1997 ,
         \pipeline/csr/N1996 , \pipeline/csr/N1995 , \pipeline/csr/N1994 ,
         \pipeline/csr/N1993 , \pipeline/csr/N1992 , \pipeline/csr/N1991 ,
         \pipeline/csr/N1990 , \pipeline/csr/N1989 , \pipeline/csr/N1988 ,
         \pipeline/csr/N1987 , \pipeline/csr/N1986 , \pipeline/csr/N1985 ,
         \pipeline/csr/N1984 , \pipeline/csr/N1983 , \pipeline/csr/N1982 ,
         \pipeline/csr/N1981 , \pipeline/csr/N1980 , \pipeline/csr/N1979 ,
         \pipeline/csr/N1978 , \pipeline/csr/N1977 , \pipeline/csr/N1976 ,
         \pipeline/csr/N1975 , \pipeline/csr/N1974 , \pipeline/csr/N1973 ,
         \pipeline/csr/N1972 , \pipeline/csr/N1971 , \pipeline/csr/N1970 ,
         \pipeline/csr/N1969 , \pipeline/csr/N1968 , \pipeline/csr/N1967 ,
         \pipeline/csr/N1966 , \pipeline/csr/N1965 , \pipeline/csr/N1964 ,
         \pipeline/csr/N1963 , \pipeline/csr/N1962 , \pipeline/csr/N1961 ,
         \pipeline/csr/N1960 , \pipeline/csr/N1959 , \pipeline/csr/N1958 ,
         \pipeline/csr/N1957 , \pipeline/csr/N1956 , \pipeline/csr/N1955 ,
         \pipeline/csr/N1954 , \pipeline/csr/N1953 , \pipeline/csr/N1952 ,
         \pipeline/csr/N1951 , \pipeline/csr/N1950 , \pipeline/csr/N1949 ,
         \pipeline/csr/N1948 , \pipeline/csr/N1947 , \pipeline/csr/N1946 ,
         \pipeline/csr/N1945 , \pipeline/csr/N1944 , \pipeline/csr/N1943 ,
         \pipeline/csr/N1942 , \pipeline/csr/N1941 , \pipeline/csr/N1940 ,
         \pipeline/csr/N1939 , \pipeline/csr/N1938 , \pipeline/csr/N1937 ,
         \pipeline/csr/N1936 , \pipeline/csr/N1935 , \pipeline/csr/N1934 ,
         \pipeline/csr/N1933 , \pipeline/csr/N1932 , \pipeline/csr/N1931 ,
         \pipeline/csr/N1930 , \pipeline/csr/N1929 , \pipeline/csr/N1928 ,
         \pipeline/csr/N1927 , \pipeline/csr/N1926 , \pipeline/csr/N1925 ,
         \pipeline/csr/N1924 , \pipeline/csr/N1923 , \pipeline/csr/N1922 ,
         \pipeline/csr/N1921 , \pipeline/csr/N1920 , \pipeline/csr/N1919 ,
         \pipeline/csr/N1918 , \pipeline/csr/N1917 , \pipeline/csr/N1916 ,
         \pipeline/csr/N1915 , \pipeline/csr/N1914 , \pipeline/csr/N1913 ,
         \pipeline/csr/N1912 , \pipeline/csr/N1911 , \pipeline/csr/N1910 ,
         \pipeline/csr/N1909 , \pipeline/csr/N1908 , \pipeline/csr/N1907 ,
         \pipeline/csr/N1906 , \pipeline/csr/N1905 , \pipeline/csr/N1904 ,
         \pipeline/csr/N1903 , \pipeline/csr/N1902 , \pipeline/csr/N1901 ,
         \pipeline/csr/N1900 , \pipeline/csr/N1899 , \pipeline/csr/N1898 ,
         \pipeline/csr/N1897 , \pipeline/csr/N1896 , \pipeline/csr/N1895 ,
         \pipeline/csr/N1894 , \pipeline/csr/N1893 , \pipeline/csr/N1892 ,
         \pipeline/csr/N1891 , \pipeline/csr/N1890 , \pipeline/csr/N1889 ,
         \pipeline/csr/N1888 , \pipeline/csr/N1887 , \pipeline/csr/N1886 ,
         \pipeline/csr/N1885 , \pipeline/csr/N1884 , \pipeline/csr/N1883 ,
         \pipeline/csr/N1882 , \pipeline/csr/N1881 , \pipeline/csr/N1880 ,
         \pipeline/csr/N1879 , \pipeline/csr/N1878 , \pipeline/csr/N1877 ,
         \pipeline/csr/N1876 , \pipeline/csr/N1875 , \pipeline/csr/N1874 ,
         \pipeline/csr/N1873 , \pipeline/csr/mcause[31] , \pipeline/csr/mip_3 ,
         \pipeline/csr/mip[7] , \pipeline/csr/system_wen ,
         \pipeline/csr/priv_stack_0 , n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8380, n8382,
         n8384, n8385, n8386, n8387, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8400, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8861, n8862,
         n8864, n8865, n8866, n8867, n8868, n8869, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10128, n10129, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10142, n10143, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
         n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
         n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
         n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
         n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
         n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
         n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
         n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
         n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
         n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
         n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
         n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
         n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
         n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,
         n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
         n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636,
         n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
         n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
         n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,
         n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
         n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676,
         n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684,
         n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
         n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,
         n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,
         n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
         n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
         n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732,
         n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
         n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748,
         n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756,
         n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,
         n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,
         n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780,
         n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788,
         n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796,
         n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804,
         n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812,
         n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820,
         n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828,
         n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836,
         n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844,
         n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852,
         n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860,
         n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868,
         n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876,
         n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884,
         n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892,
         n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900,
         n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908,
         n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916,
         n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924,
         n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932,
         n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940,
         n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948,
         n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956,
         n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964,
         n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972,
         n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980,
         n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,
         n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996,
         n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,
         n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012,
         n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020,
         n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028,
         n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036,
         n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044,
         n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052,
         n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060,
         n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068,
         n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,
         n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084,
         n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092,
         n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100,
         n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108,
         n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116,
         n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124,
         n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132,
         n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140,
         n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,
         n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156,
         n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164,
         n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172,
         n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180,
         n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188,
         n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196,
         n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204,
         n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212,
         n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220,
         n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228,
         n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236,
         n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244,
         n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252,
         n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260,
         n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268,
         n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276,
         n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284,
         n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
         n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300,
         n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308,
         n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316,
         n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324,
         n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332,
         n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340,
         n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348,
         n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356,
         n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364,
         n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372,
         n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380,
         n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388,
         n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396,
         n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404,
         n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412,
         n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420,
         n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428,
         n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436,
         n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444,
         n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452,
         n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460,
         n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468,
         n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476,
         n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484,
         n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492,
         n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500,
         n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508,
         n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516,
         n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524,
         n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532,
         n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540,
         n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548,
         n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556,
         n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564,
         n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572,
         n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580,
         n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588,
         n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596,
         n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604,
         n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612,
         n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620,
         n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628,
         n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636,
         n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644,
         n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652,
         n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660,
         n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668,
         n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
         n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684,
         n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692,
         n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700,
         n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708,
         n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716,
         n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724,
         n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732,
         n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740,
         n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748,
         n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756,
         n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764,
         n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772,
         n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780,
         n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788,
         n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796,
         n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804,
         n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812,
         n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820,
         n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828,
         n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836,
         n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844,
         n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852,
         n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860,
         n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868,
         n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876,
         n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884,
         n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892,
         n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900,
         n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908,
         n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916,
         n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924,
         n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932,
         n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940,
         n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948,
         n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956,
         n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964,
         n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972,
         n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980,
         n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988,
         n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996,
         n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004,
         n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012,
         n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020,
         n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028,
         n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036,
         n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044,
         n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052,
         n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060,
         n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068,
         n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076,
         n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084,
         n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092,
         n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100,
         n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108,
         n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116,
         n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124,
         n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132,
         n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140,
         n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148,
         n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156,
         n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164,
         n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172,
         n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180,
         n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188,
         n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196,
         n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204,
         n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212,
         n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220,
         n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228,
         n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236,
         n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244,
         n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252,
         n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260,
         n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268,
         n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276,
         n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284,
         n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292,
         n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300,
         n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308,
         n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316,
         n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324,
         n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332,
         n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340,
         n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348,
         n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356,
         n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364,
         n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372,
         n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380,
         n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388,
         n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396,
         n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404,
         n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412,
         n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420,
         n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428,
         n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436,
         n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444,
         n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452,
         n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460,
         n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468,
         n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476,
         n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484,
         n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492,
         n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500,
         n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508,
         n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516,
         n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524,
         n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532,
         n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540,
         n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548,
         n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556,
         n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564,
         n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572,
         n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580,
         n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588,
         n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596,
         n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604,
         n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612,
         n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620,
         n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628,
         n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636,
         n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644,
         n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652,
         n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660,
         n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668,
         n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676,
         n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684,
         n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692,
         n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700,
         n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708,
         n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716,
         n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724,
         n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732,
         n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740,
         n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748,
         n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756,
         n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764,
         n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772,
         n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780,
         n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788,
         n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796,
         n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804,
         n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812,
         n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820,
         n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828,
         n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836,
         n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844,
         n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852,
         n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860,
         n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868,
         n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876,
         n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884,
         n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892,
         n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900,
         n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908,
         n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916,
         n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924,
         n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932,
         n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940,
         n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948,
         n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956,
         n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964,
         n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972,
         n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980,
         n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988,
         n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996,
         n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004,
         n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012,
         n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020,
         n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028,
         n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036,
         n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044,
         n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052,
         n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060,
         n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068,
         n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076,
         n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084,
         n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092,
         n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100,
         n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108,
         n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116,
         n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124,
         n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132,
         n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140,
         n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148,
         n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156,
         n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164,
         n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172,
         n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180,
         n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188,
         n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196,
         n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204,
         n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212,
         n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220,
         n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228,
         n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236,
         n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244,
         n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252,
         n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260,
         n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268,
         n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276,
         n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284,
         n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292,
         n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300,
         n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308,
         n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316,
         n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324,
         n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332,
         n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340,
         n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348,
         n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356,
         n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364,
         n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372,
         n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380,
         n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388,
         n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396,
         n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404,
         n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412,
         n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420,
         n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428,
         n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436,
         n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444,
         n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452,
         n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460,
         n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468,
         n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476,
         n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484,
         n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492,
         n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500,
         n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508,
         n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516,
         n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524,
         n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532,
         n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540,
         n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548,
         n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556,
         n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564,
         n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572,
         n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580,
         n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588,
         n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596,
         n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604,
         n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612,
         n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620,
         n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628,
         n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636,
         n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644,
         n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652,
         n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660,
         n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668,
         n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676,
         n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684,
         n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692,
         n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700,
         n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708,
         n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716,
         n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724,
         n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732,
         n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740,
         n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748,
         n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756,
         n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764,
         n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772,
         n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780,
         n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788,
         n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796,
         n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804,
         n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812,
         n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820,
         n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828,
         n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836,
         n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844,
         n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852,
         n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860,
         n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868,
         n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876,
         n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884,
         n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892,
         n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900,
         n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908,
         n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916,
         n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924,
         n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932,
         n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940,
         n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948,
         n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956,
         n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964,
         n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972,
         n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980,
         n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988,
         n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996,
         n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004,
         n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012,
         n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020,
         n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028,
         n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036,
         n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044,
         n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052,
         n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060,
         n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068,
         n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076,
         n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084,
         n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092,
         n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100,
         n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108,
         n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116,
         n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124,
         n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132,
         n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140,
         n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148,
         n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156,
         n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164,
         n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172,
         n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180,
         n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188,
         n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196,
         n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204,
         n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212,
         n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220,
         n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228,
         n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236,
         n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244,
         n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252,
         n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260,
         n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268,
         n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276,
         n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284,
         n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292,
         n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300,
         n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308,
         n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316,
         n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324,
         n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332,
         n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340,
         n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348,
         n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356,
         n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364,
         n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372,
         n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380,
         n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388,
         n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396,
         n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404,
         n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412,
         n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420,
         n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428,
         n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436,
         n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444,
         n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452,
         n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460,
         n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468,
         n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476,
         n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484,
         n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492,
         n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500,
         n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508,
         n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516,
         n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524,
         n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532,
         n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540,
         n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548,
         n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556,
         n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564,
         n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572,
         n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580,
         n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588,
         n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596,
         n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604,
         n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612,
         n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620,
         n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628,
         n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636,
         n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644,
         n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652,
         n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660,
         n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668,
         n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676,
         n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684,
         n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692,
         n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700,
         n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708,
         n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716,
         n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724,
         n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732,
         n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740,
         n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748,
         n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756,
         n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764,
         n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772,
         n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780,
         n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788,
         n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796,
         n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804,
         n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812,
         n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820,
         n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828,
         n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836,
         n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844,
         n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852,
         n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860,
         n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868,
         n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876,
         n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884,
         n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892,
         n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900,
         n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908,
         n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916,
         n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924,
         n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932,
         n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940,
         n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948,
         n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956,
         n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964,
         n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972,
         n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980,
         n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988,
         n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996,
         n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004,
         n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012,
         n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020,
         n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028,
         n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036,
         n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044,
         n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052,
         n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060,
         n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068,
         n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076,
         n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084,
         n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092,
         n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100,
         n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108,
         n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116,
         n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124,
         n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132,
         n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140,
         n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148,
         n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156,
         n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164,
         n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172,
         n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180,
         n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188,
         n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196,
         n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204,
         n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212,
         n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220,
         n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228,
         n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236,
         n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244,
         n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252,
         n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260,
         n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268,
         n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276,
         n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284,
         n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292,
         n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300,
         n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308,
         n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316,
         n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324,
         n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332,
         n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340,
         n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348,
         n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356,
         n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364,
         n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372,
         n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380,
         n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388,
         n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396,
         n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404,
         n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412,
         n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420,
         n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428,
         n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436,
         n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444,
         n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452,
         n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460,
         n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468,
         n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476,
         n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484,
         n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492,
         n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500,
         n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508,
         n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516,
         n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524,
         n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532,
         n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540,
         n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548,
         n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556,
         n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564,
         n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572,
         n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580,
         n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588,
         n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596,
         n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604,
         n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612,
         n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620,
         n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628,
         n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636,
         n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644,
         n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652,
         n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660,
         n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668,
         n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676,
         n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684,
         n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692,
         n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700,
         n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708,
         n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716,
         n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724,
         n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732,
         n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740,
         n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748,
         n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756,
         n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764,
         n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772,
         n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780,
         n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788,
         n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796,
         n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804,
         n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812,
         n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820,
         n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828,
         n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836,
         n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844,
         n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852,
         n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860,
         n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868,
         n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876,
         n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884,
         n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892,
         n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900,
         n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908,
         n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916,
         n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924,
         n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932,
         n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940,
         n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948,
         n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956,
         n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964,
         n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972,
         n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980,
         n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988,
         n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996,
         n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004,
         n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012,
         n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020,
         n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028,
         n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036,
         n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044,
         n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052,
         n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060,
         n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068,
         n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076,
         n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084,
         n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092,
         n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100,
         n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108,
         n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116,
         n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124,
         n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132,
         n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140,
         n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148,
         n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156,
         n21157, n21158, n21159, n21160, n21161, n21162, n21163, n21164,
         n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172,
         n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180,
         n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188,
         n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196,
         n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204,
         n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212,
         n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220,
         n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228,
         n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236,
         n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244,
         n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252,
         n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260,
         n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268,
         n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276,
         n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284,
         n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292,
         n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300,
         n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308,
         n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316,
         n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324,
         n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332,
         n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340,
         n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348,
         n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356,
         n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364,
         n21365, n21366, n21367, n21368, n21369, n21370, n21371, n21372,
         n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380,
         n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388,
         n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21396,
         n21397, n21398, n21399, n21400, n21401, n21402, n21403, n21404,
         n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412,
         n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420,
         n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428,
         n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436,
         n21437, n21438, n21439, n21440, n21441, n21442, n21443, n21444,
         n21445, n21446, n21447, n21448, n21449, n21450, n21451, n21452,
         n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460,
         n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468,
         n21469, n21470, n21471, n21472, n21473, n21474, n21475, n21476,
         n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484,
         n21485, n21486, n21487, n21488, n21489, n21490, n21491, n21492,
         n21493, n21494, n21495, n21496, n21497, n21498, n21499, n21500,
         n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508,
         n21509, n21510, n21511, n21512, n21513, n21514, n21515, n21516,
         n21517, n21518, n21519, n21520, n21521, n21522, n21523, n21524,
         n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532,
         n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540,
         n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548,
         n21549, n21550, n21551, n21552, n21553, n21554, n21555, n21556,
         n21557, n21558, n21559, n21560, n21561, n21562, n21563, n21564,
         n21565, n21566, n21567, n21568, n21569, n21570, n21571, n21572,
         n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580,
         n21581, n21582, n21583, n21584, n21585, n21586, n21587, n21588,
         n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596,
         n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604,
         n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612,
         n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620,
         n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628,
         n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636,
         n21637, n21638, n21639, n21640, n21641, n21642, n21643, n21644,
         n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652,
         n21653, n21654, n21655, n21656, n21657, n21658, n21659, n21660,
         n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21668,
         n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676,
         n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684,
         n21685, n21686, n21687, n21688, n21689, n21690, n21691, n21692,
         n21693, n21694, n21695, n21696, n21697, n21698, n21699, n21700,
         n21701, n21702, n21703, n21704, n21705, n21706, n21707, n21708,
         n21709, n21710, n21711, n21712, n21713, n21714, n21715, n21716,
         n21717, n21718, n21719, n21720, n21721, n21722, n21723, n21724,
         n21725, n21726, n21727, n21728, n21729, n21730, n21731, n21732,
         n21733, n21734, n21735, n21736, n21737, n21738, n21739, n21740,
         n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748,
         n21749, n21750, n21751, n21752, n21753, n21754, n21755, n21756,
         n21757, n21758, n21759, n21760, n21761, n21762, n21763, n21764,
         n21765, n21766, n21767, n21768, n21769, n21770, n21771, n21772,
         n21773, n21774, n21775, n21776, n21777, n21778, n21779, n21780,
         n21781, n21782, n21783, n21784, n21785, n21786, n21787, n21788,
         n21789, n21790, n21791, n21792, n21793, n21794, n21795, n21796,
         n21797, n21798, n21799, n21800, n21801, n21802, n21803, n21804,
         n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812,
         n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820,
         n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828,
         n21829, n21830, n21831, n21832, n21833, n21834, n21835, n21836,
         n21837, n21838, n21839, n21840, n21841, n21842, n21843, n21844,
         n21845, n21846, n21847, n21848, n21849, n21850, n21851, n21852,
         n21853, n21854, n21855, n21856, n21857, n21858, n21859, n21860,
         n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868,
         n21869, n21870, n21871, n21872, n21873, n21874, n21875, n21876,
         n21877, n21878, n21879, n21880, n21881, n21882, n21883, n21884,
         n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892,
         n21893, n21894, n21895, n21896, n21897, n21898, n21899, n21900,
         n21901, n21902, n21903, n21904, n21905, n21906, n21907, n21908,
         n21909, n21910, n21911, n21912, n21913, n21914, n21915, n21916,
         n21917, n21918, n21919, n21920, n21921, n21922, n21923, n21924,
         n21925, n21926, n21927, n21928, n21929, n21930, n21931, n21932,
         n21933, n21934, n21935, n21936, n21937, n21938, n21939, n21940,
         n21941, n21942, n21943, n21944, n21945, n21946, n21947, n21948,
         n21949, n21950, n21951, n21952, n21953, n21954, n21955, n21956,
         n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964,
         n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972,
         n21973, n21974, n21975, n21976, n21977, n21978, n21979, n21980,
         n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988,
         n21989, n21990, n21991, n21992, n21993, n21994, n21995, n21996,
         n21997, n21998, n21999, n22000, n22001, n22002, n22003, n22004,
         n22005, n22006, n22007, n22008, n22009, n22010, n22011, n22012,
         n22013, n22014, n22015, n22016, n22017, n22018, n22019, n22020,
         n22021, n22022, n22023, n22024, n22025, n22026, n22027, n22028,
         n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036,
         n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044,
         n22045, n22046, n22047, n22048, n22049, n22050, n22051, n22052,
         n22053, n22054, n22055, n22056, n22057, n22058, n22059, n22060,
         n22061, n22062, n22063, n22064, n22065, n22066, n22067, n22068,
         n22069, n22070, n22071, n22072, n22073, n22074, n22075, n22076,
         n22077, n22078, n22079, n22080, n22081, n22082, n22083, n22084,
         n22085, n22086, n22087, n22088, n22089, n22090, n22091, n22092,
         n22093, n22094, n22095, n22096, n22097, n22098, n22099, n22100,
         n22101, n22102, n22103, n22104, n22105, n22106, n22107, n22108,
         n22109, n22110, n22111, n22112, n22113, n22114, n22115, n22116,
         n22117, n22118, n22119, n22120, n22121, n22122, n22123, n22124,
         n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132,
         n22133, n22134, n22135, n22136, n22137, n22138, n22139, n22140,
         n22141, n22142, n22143, n22144, n22145, n22146, n22147, n22148,
         n22149, n22150, n22151, n22152, n22153, n22154, n22155, n22156,
         n22157, n22158, n22159, n22160, n22161, n22162, n22163, n22164,
         n22165, n22166, n22167, n22168, n22169, n22170, n22171, n22172,
         n22173, n22174, n22175, n22176, n22177, n22178, n22179, n22180,
         n22181, n22182, n22183, n22184, n22185, n22186, n22187, n22188,
         n22189, n22190, n22191, n22192, n22193, n22194, n22195, n22196,
         n22197, n22198, n22199, n22200, n22201, n22202, n22203, n22204,
         n22205, n22206, n22207, n22208, n22209, n22210, n22211, n22212,
         n22213, n22214, n22215, n22216, n22217, n22218, n22219, n22220,
         n22221, n22222, n22223, n22224, n22225, n22226, n22227, n22228,
         n22229, n22230, n22231, n22232, n22233, n22234, n22235, n22236,
         n22237, n22238, n22239, n22240, n22241, n22242, n22243, n22244,
         n22245, n22246, n22247, n22248, n22249, n22250, n22251, n22252,
         n22253, n22254, n22255, n22256, n22257, n22258, n22259, n22260,
         n22261, n22262, n22263, n22264, n22265, n22266, n22267, n22268,
         n22269, n22270, n22271, n22272, n22273, n22274, n22275, n22276,
         n22277, n22278, n22279, n22280, n22281, n22282, n22283, n22284,
         n22285, n22286, n22287, n22288, n22289, n22290, n22291, n22292,
         n22293, n22294, n22295, n22296, n22297, n22298, n22299, n22300,
         n22301, n22302, n22303, n22304, n22305, n22306, n22307, n22308,
         n22309, n22310, n22311, n22312, n22313, n22314, n22315, n22316,
         n22317, n22318, n22319, n22320, n22321, n22322, n22323, n22324,
         n22325, n22326, n22327, n22328, n22329, n22330, n22331, n22332,
         n22333, n22334, n22335, n22336, n22337, n22338, n22339, n22340,
         n22341, n22342, n22343, n22344, n22345, n22346, n22347, n22348,
         n22349, n22350, n22351, n22352, n22353, n22354, n22355, n22356,
         n22357, n22358, n22359, n22360, n22361, n22362, n22363, n22364,
         n22365, n22366, n22367, n22368, n22369, n22370, n22371, n22372,
         n22373, n22374, n22375, n22376, n22377, n22378, n22379, n22380,
         n22381, n22382, n22383, n22384, n22385, n22386, n22387, n22388,
         n22389, n22390, n22391, n22392, n22393, n22394, n22395, n22396,
         n22397, n22398, n22399, n22400, n22401, n22402, n22403, n22404,
         n22405, n22406, n22407, n22408, n22409, n22410, n22411, n22412,
         n22413, n22414, n22415, n22416, n22417, n22418, n22419, n22420,
         n22421, n22422, n22423, n22424, n22425, n22426, n22427, n22428,
         n22429, n22430, n22431, n22432, n22433, n22434, n22435, n22436,
         n22437, n22438, n22439, n22440, n22441, n22442, n22443, n22444,
         n22445, n22446, n22447, n22448, n22449, n22450, n22451, n22452,
         n22453, n22454, n22455, n22456, n22457, n22458, n22459, n22460,
         n22461, n22462, n22463, n22464, n22465, n22466, n22467, n22468,
         n22469, n22470, n22471, n22472, n22473, n22474, n22475, n22476,
         n22477, n22478, n22479, n22480, n22481, n22482, n22483, n22484,
         n22485, n22486, n22487, n22488, n22489, n22490, n22491, n22492,
         n22493, n22494, n22495, n22496, n22497, n22498, n22499, n22500,
         n22501, n22502, n22503, n22504, n22505, n22506, n22507, n22508,
         n22509, n22510, n22511, n22512, n22513, n22514, n22515, n22516,
         n22517, n22518, n22519, n22520, n22521, n22522, n22523, n22524,
         n22525, n22526, n22527, n22528, n22529, n22530, n22531, n22532,
         n22533, n22534, n22535, n22536, n22537, n22538, n22539, n22540,
         n22541, n22542, n22543, n22544, n22545, n22546, n22547, n22548,
         n22549, n22550, n22551, n22552, n22553, n22554, n22555, n22556,
         n22557, n22558, n22559, n22560, n22561, n22562, n22563, n22564,
         n22565, n22566, n22567, n22568, n22569, n22570, n22571, n22572,
         n22573, n22574, n22575, n22576, n22577, n22578, n22579, n22580,
         n22581, n22582, n22583, n22584, n22585, n22586, n22587, n22588,
         n22589, n22590, n22591, n22592, n22593, n22594, n22595, n22596,
         n22597, n22598, n22599, n22600, n22601, n22602, n22603, n22604,
         n22605, n22606, n22607, n22608, n22609, n22610, n22611, n22612,
         n22613, n22614, n22615, n22616, n22617, n22618, n22619, n22620,
         n22621, n22622, n22623, n22624, n22625, n22626, n22627, n22628,
         n22629, n22630, n22631, n22632, n22633, n22634, n22635, n22636,
         n22637, n22638, n22639, n22640, n22641, n22642, n22643, n22644,
         n22645, n22646, n22647, n22648, n22649, n22650, n22651, n22652,
         n22653, n22654, n22655, n22656, n22657, n22658, n22659, n22660,
         n22661, n22662, n22663, n22664, n22665, n22666, n22667, n22668,
         n22669, n22670, n22671, n22672, n22673, n22674, n22675, n22676,
         n22677, n22678, n22679, n22680, n22681, n22682, n22683, n22684,
         n22685, n22686, n22687, n22688, n22689, n22690, n22691, n22692,
         n22693, n22694, n22695, n22696, n22697, n22698, n22699, n22700,
         n22701, n22702, n22703, n22704, n22705, n22706, n22707, n22708,
         n22709, n22710, n22711, n22712, n22713, n22714, n22715, n22716,
         n22717, n22718, n22719, n22720, n22721, n22722, n22723, n22724,
         n22725, n22726, n22727, n22728, n22729, n22730, n22731, n22732,
         n22733, n22734, n22735, n22736, n22737, n22738, n22739, n22740,
         n22741, n22742, n22743, n22744, n22745, n22746, n22747, n22748,
         n22749, n22750, n22751, n22752, n22753, n22754, n22755, n22756,
         n22757, n22758, n22759, n22850, n22851, n22852, n22853, n22854,
         n22855, n22856, n22857, n22858, n22859, n22860, n22861, n22862,
         n22863, n22866, n22896, n22898;
  wire   [31:0] imem_rdata;
  wire   [31:0] dmem_rdata;
  wire   [2:0] \pipeline/dmem_type_WB ;
  wire   [31:0] \pipeline/csr_rdata_WB ;
  wire   [31:0] \pipeline/alu_out_WB ;
  wire   [31:8] \pipeline/store_data_WB ;
  wire   [31:0] \pipeline/PC_WB ;
  wire   [31:0] \pipeline/md_resp_result ;
  wire   [31:0] \pipeline/epc ;
  wire   [31:0] \pipeline/PC_DX ;
  wire   [31:0] \pipeline/PC_IF ;
  wire   [1:0] \pipeline/prv ;
  wire   [1:0] \pipeline/wb_src_sel_WB ;
  wire   [4:0] \pipeline/reg_to_wr_WB ;
  wire   [31:0] \pipeline/inst_DX ;
  wire   [3:0] \pipeline/ctrl/prev_ex_code_WB ;
  wire   [1:0] \pipeline/md/op ;
  wire   [4:0] \pipeline/md/counter ;
  wire   [1:0] \pipeline/md/out_sel ;
  wire   [63:0] \pipeline/md/b ;
  wire   [63:0] \pipeline/md/a ;
  wire   [63:32] \pipeline/md/result ;
  wire   [1:0] \pipeline/md/state ;
  wire   [31:0] \pipeline/csr/mscratch ;
  wire   [63:0] \pipeline/csr/instret_full ;
  wire   [63:0] \pipeline/csr/time_full ;
  wire   [63:0] \pipeline/csr/cycle_full ;
  wire   [31:0] \pipeline/csr/from_host ;
  wire   [31:0] \pipeline/csr/to_host ;
  wire   [31:0] \pipeline/csr/mbadaddr ;
  wire   [3:0] \pipeline/csr/mecode ;
  wire   [63:0] \pipeline/csr/mtime_full ;
  wire   [31:0] \pipeline/csr/mtimecmp ;
  wire   [31:0] \pipeline/csr/mie ;
  wire   [5:3] \pipeline/csr/priv_stack ;
  wire   [31:0] \pipeline/csr/mtvec ;
  assign htif_debug_stats_pcr = 1'b0;
  assign htif_pcr_resp_data[63] = 1'b0;
  assign imem_rdata[31] = imem_hrdata[31];
  assign imem_rdata[30] = imem_hrdata[30];
  assign imem_rdata[29] = imem_hrdata[29];
  assign imem_rdata[28] = imem_hrdata[28];
  assign imem_rdata[27] = imem_hrdata[27];
  assign imem_rdata[26] = imem_hrdata[26];
  assign imem_rdata[25] = imem_hrdata[25];
  assign imem_rdata[24] = imem_hrdata[24];
  assign imem_rdata[23] = imem_hrdata[23];
  assign imem_rdata[22] = imem_hrdata[22];
  assign imem_rdata[21] = imem_hrdata[21];
  assign imem_rdata[20] = imem_hrdata[20];
  assign imem_rdata[19] = imem_hrdata[19];
  assign imem_rdata[18] = imem_hrdata[18];
  assign imem_rdata[17] = imem_hrdata[17];
  assign imem_rdata[16] = imem_hrdata[16];
  assign imem_rdata[15] = imem_hrdata[15];
  assign imem_rdata[14] = imem_hrdata[14];
  assign imem_rdata[13] = imem_hrdata[13];
  assign imem_rdata[12] = imem_hrdata[12];
  assign imem_rdata[11] = imem_hrdata[11];
  assign imem_rdata[10] = imem_hrdata[10];
  assign imem_rdata[9] = imem_hrdata[9];
  assign imem_rdata[8] = imem_hrdata[8];
  assign imem_rdata[7] = imem_hrdata[7];
  assign imem_rdata[6] = imem_hrdata[6];
  assign imem_rdata[5] = imem_hrdata[5];
  assign imem_rdata[4] = imem_hrdata[4];
  assign imem_rdata[3] = imem_hrdata[3];
  assign imem_rdata[2] = imem_hrdata[2];
  assign imem_rdata[1] = imem_hrdata[1];
  assign imem_rdata[0] = imem_hrdata[0];
  assign imem_badmem_e = imem_hresp[0];
  assign dmem_rdata[31] = dmem_hrdata[31];
  assign dmem_rdata[30] = dmem_hrdata[30];
  assign dmem_rdata[29] = dmem_hrdata[29];
  assign dmem_rdata[28] = dmem_hrdata[28];
  assign dmem_rdata[27] = dmem_hrdata[27];
  assign dmem_rdata[26] = dmem_hrdata[26];
  assign dmem_rdata[25] = dmem_hrdata[25];
  assign dmem_rdata[24] = dmem_hrdata[24];
  assign dmem_rdata[23] = dmem_hrdata[23];
  assign dmem_rdata[22] = dmem_hrdata[22];
  assign dmem_rdata[21] = dmem_hrdata[21];
  assign dmem_rdata[20] = dmem_hrdata[20];
  assign dmem_rdata[19] = dmem_hrdata[19];
  assign dmem_rdata[18] = dmem_hrdata[18];
  assign dmem_rdata[17] = dmem_hrdata[17];
  assign dmem_rdata[16] = dmem_hrdata[16];
  assign dmem_rdata[15] = dmem_hrdata[15];
  assign dmem_rdata[14] = dmem_hrdata[14];
  assign dmem_rdata[13] = dmem_hrdata[13];
  assign dmem_rdata[12] = dmem_hrdata[12];
  assign dmem_rdata[11] = dmem_hrdata[11];
  assign dmem_rdata[10] = dmem_hrdata[10];
  assign dmem_rdata[9] = dmem_hrdata[9];
  assign dmem_rdata[8] = dmem_hrdata[8];
  assign dmem_rdata[7] = dmem_hrdata[7];
  assign dmem_rdata[6] = dmem_hrdata[6];
  assign dmem_rdata[5] = dmem_hrdata[5];
  assign dmem_rdata[4] = dmem_hrdata[4];
  assign dmem_rdata[3] = dmem_hrdata[3];
  assign dmem_rdata[2] = dmem_hrdata[2];
  assign dmem_rdata[1] = dmem_hrdata[1];
  assign dmem_rdata[0] = dmem_hrdata[0];
  assign dmem_badmem_e = dmem_hresp[0];
  assign htif_ipi_resp_ready = 1'b1;
  assign htif_ipi_req_data = 1'b0;
  assign htif_ipi_req_valid = 1'b0;
  assign htif_pcr_resp_data[32] = 1'b0;
  assign htif_pcr_resp_data[33] = 1'b0;
  assign htif_pcr_resp_data[34] = 1'b0;
  assign htif_pcr_resp_data[35] = 1'b0;
  assign htif_pcr_resp_data[36] = 1'b0;
  assign htif_pcr_resp_data[37] = 1'b0;
  assign htif_pcr_resp_data[38] = 1'b0;
  assign htif_pcr_resp_data[39] = 1'b0;
  assign htif_pcr_resp_data[40] = 1'b0;
  assign htif_pcr_resp_data[41] = 1'b0;
  assign htif_pcr_resp_data[42] = 1'b0;
  assign htif_pcr_resp_data[43] = 1'b0;
  assign htif_pcr_resp_data[44] = 1'b0;
  assign htif_pcr_resp_data[45] = 1'b0;
  assign htif_pcr_resp_data[46] = 1'b0;
  assign htif_pcr_resp_data[47] = 1'b0;
  assign htif_pcr_resp_data[48] = 1'b0;
  assign htif_pcr_resp_data[49] = 1'b0;
  assign htif_pcr_resp_data[50] = 1'b0;
  assign htif_pcr_resp_data[51] = 1'b0;
  assign htif_pcr_resp_data[52] = 1'b0;
  assign htif_pcr_resp_data[53] = 1'b0;
  assign htif_pcr_resp_data[54] = 1'b0;
  assign htif_pcr_resp_data[55] = 1'b0;
  assign htif_pcr_resp_data[56] = 1'b0;
  assign htif_pcr_resp_data[57] = 1'b0;
  assign htif_pcr_resp_data[58] = 1'b0;
  assign htif_pcr_resp_data[59] = 1'b0;
  assign htif_pcr_resp_data[60] = 1'b0;
  assign htif_pcr_resp_data[61] = 1'b0;
  assign htif_pcr_resp_data[62] = 1'b0;
  assign dmem_htrans[0] = 1'b0;
  assign dmem_hprot[0] = 1'b0;
  assign dmem_hprot[1] = 1'b0;
  assign dmem_hprot[2] = 1'b0;
  assign dmem_hprot[3] = 1'b0;
  assign dmem_hmastlock = 1'b0;
  assign dmem_hburst[0] = 1'b0;
  assign dmem_hburst[1] = 1'b0;
  assign dmem_hburst[2] = 1'b0;
  assign dmem_hsize[2] = 1'b0;
  assign imem_hwdata[0] = 1'b0;
  assign imem_hwdata[1] = 1'b0;
  assign imem_hwdata[2] = 1'b0;
  assign imem_hwdata[3] = 1'b0;
  assign imem_hwdata[4] = 1'b0;
  assign imem_hwdata[5] = 1'b0;
  assign imem_hwdata[6] = 1'b0;
  assign imem_hwdata[7] = 1'b0;
  assign imem_hwdata[8] = 1'b0;
  assign imem_hwdata[9] = 1'b0;
  assign imem_hwdata[10] = 1'b0;
  assign imem_hwdata[11] = 1'b0;
  assign imem_hwdata[12] = 1'b0;
  assign imem_hwdata[13] = 1'b0;
  assign imem_hwdata[14] = 1'b0;
  assign imem_hwdata[15] = 1'b0;
  assign imem_hwdata[16] = 1'b0;
  assign imem_hwdata[17] = 1'b0;
  assign imem_hwdata[18] = 1'b0;
  assign imem_hwdata[19] = 1'b0;
  assign imem_hwdata[20] = 1'b0;
  assign imem_hwdata[21] = 1'b0;
  assign imem_hwdata[22] = 1'b0;
  assign imem_hwdata[23] = 1'b0;
  assign imem_hwdata[24] = 1'b0;
  assign imem_hwdata[25] = 1'b0;
  assign imem_hwdata[26] = 1'b0;
  assign imem_hwdata[27] = 1'b0;
  assign imem_hwdata[28] = 1'b0;
  assign imem_hwdata[29] = 1'b0;
  assign imem_hwdata[30] = 1'b0;
  assign imem_hwdata[31] = 1'b0;
  assign imem_htrans[0] = 1'b0;
  assign imem_htrans[1] = 1'b1;
  assign imem_hprot[0] = 1'b0;
  assign imem_hprot[1] = 1'b0;
  assign imem_hprot[2] = 1'b0;
  assign imem_hprot[3] = 1'b0;
  assign imem_hmastlock = 1'b0;
  assign imem_hburst[0] = 1'b0;
  assign imem_hburst[1] = 1'b0;
  assign imem_hburst[2] = 1'b0;
  assign imem_hsize[0] = 1'b0;
  assign imem_hsize[1] = 1'b1;
  assign imem_hsize[2] = 1'b0;
  assign imem_hwrite = 1'b0;

  or2_1 \pipeline/csr/C4919  ( .ip1(n22898), .ip2(n22896), .op(
        \pipeline/csr/system_wen ) );
  and2_1 \pipeline/csr/C4923  ( .ip1(n22866), .ip2(n10143), .op(
        \pipeline/csr/N2385 ) );
  and2_1 \pipeline/csr/C4925  ( .ip1(n22866), .ip2(n10142), .op(
        \pipeline/csr/N2387 ) );
  dp_1 \pipeline/md/result_reg[0]  ( .ip(n8634), .ck(clk), .q(
        \pipeline/md_resp_result [0]) );
  dp_1 \pipeline/md/result_reg[1]  ( .ip(n8633), .ck(clk), .q(
        \pipeline/md_resp_result [1]) );
  dp_1 \pipeline/md/result_reg[2]  ( .ip(n8632), .ck(clk), .q(
        \pipeline/md_resp_result [2]) );
  dp_1 \pipeline/md/result_reg[3]  ( .ip(n8631), .ck(clk), .q(
        \pipeline/md_resp_result [3]) );
  dp_1 \pipeline/md/result_reg[4]  ( .ip(n8630), .ck(clk), .q(
        \pipeline/md_resp_result [4]) );
  dp_1 \pipeline/md/result_reg[5]  ( .ip(n8629), .ck(clk), .q(
        \pipeline/md_resp_result [5]) );
  dp_1 \pipeline/md/result_reg[6]  ( .ip(n8628), .ck(clk), .q(
        \pipeline/md_resp_result [6]) );
  dp_1 \pipeline/md/result_reg[7]  ( .ip(n8627), .ck(clk), .q(
        \pipeline/md_resp_result [7]) );
  dp_1 \pipeline/md/result_reg[8]  ( .ip(n8626), .ck(clk), .q(
        \pipeline/md_resp_result [8]) );
  dp_1 \pipeline/md/result_reg[9]  ( .ip(n8625), .ck(clk), .q(
        \pipeline/md_resp_result [9]) );
  dp_1 \pipeline/md/result_reg[10]  ( .ip(n8624), .ck(clk), .q(
        \pipeline/md_resp_result [10]) );
  dp_1 \pipeline/md/result_reg[11]  ( .ip(n8623), .ck(clk), .q(
        \pipeline/md_resp_result [11]) );
  dp_1 \pipeline/md/result_reg[12]  ( .ip(n8622), .ck(clk), .q(
        \pipeline/md_resp_result [12]) );
  dp_1 \pipeline/md/result_reg[13]  ( .ip(n8621), .ck(clk), .q(
        \pipeline/md_resp_result [13]) );
  dp_1 \pipeline/md/result_reg[14]  ( .ip(n8620), .ck(clk), .q(
        \pipeline/md_resp_result [14]) );
  dp_1 \pipeline/md/result_reg[15]  ( .ip(n8619), .ck(clk), .q(
        \pipeline/md_resp_result [15]) );
  dp_1 \pipeline/md/result_reg[16]  ( .ip(n8618), .ck(clk), .q(
        \pipeline/md_resp_result [16]) );
  dp_1 \pipeline/md/result_reg[17]  ( .ip(n8617), .ck(clk), .q(
        \pipeline/md_resp_result [17]) );
  dp_1 \pipeline/md/result_reg[18]  ( .ip(n8616), .ck(clk), .q(
        \pipeline/md_resp_result [18]) );
  dp_1 \pipeline/md/result_reg[19]  ( .ip(n8615), .ck(clk), .q(
        \pipeline/md_resp_result [19]) );
  dp_1 \pipeline/md/result_reg[20]  ( .ip(n8614), .ck(clk), .q(
        \pipeline/md_resp_result [20]) );
  dp_1 \pipeline/md/result_reg[21]  ( .ip(n8613), .ck(clk), .q(
        \pipeline/md_resp_result [21]) );
  dp_1 \pipeline/md/result_reg[22]  ( .ip(n8612), .ck(clk), .q(
        \pipeline/md_resp_result [22]) );
  dp_1 \pipeline/md/result_reg[23]  ( .ip(n8611), .ck(clk), .q(
        \pipeline/md_resp_result [23]) );
  dp_1 \pipeline/md/result_reg[24]  ( .ip(n8610), .ck(clk), .q(
        \pipeline/md_resp_result [24]) );
  dp_1 \pipeline/md/result_reg[25]  ( .ip(n8609), .ck(clk), .q(
        \pipeline/md_resp_result [25]) );
  dp_1 \pipeline/md/result_reg[26]  ( .ip(n8608), .ck(clk), .q(
        \pipeline/md_resp_result [26]) );
  dp_1 \pipeline/md/result_reg[27]  ( .ip(n8607), .ck(clk), .q(
        \pipeline/md_resp_result [27]) );
  dp_1 \pipeline/md/result_reg[28]  ( .ip(n8606), .ck(clk), .q(
        \pipeline/md_resp_result [28]) );
  dp_1 \pipeline/md/result_reg[29]  ( .ip(n8605), .ck(clk), .q(
        \pipeline/md_resp_result [29]) );
  dp_1 \pipeline/md/result_reg[30]  ( .ip(n8604), .ck(clk), .q(
        \pipeline/md_resp_result [30]) );
  dp_1 \pipeline/md/result_reg[31]  ( .ip(n8603), .ck(clk), .q(
        \pipeline/md_resp_result [31]) );
  dp_1 \pipeline/md/result_reg[32]  ( .ip(n8602), .ck(clk), .q(
        \pipeline/md/result [32]) );
  dp_1 \pipeline/md/result_reg[33]  ( .ip(n8601), .ck(clk), .q(
        \pipeline/md/result [33]) );
  dp_1 \pipeline/md/result_reg[34]  ( .ip(n8600), .ck(clk), .q(
        \pipeline/md/result [34]) );
  dp_1 \pipeline/md/result_reg[35]  ( .ip(n8599), .ck(clk), .q(
        \pipeline/md/result [35]) );
  dp_1 \pipeline/md/result_reg[36]  ( .ip(n8598), .ck(clk), .q(
        \pipeline/md/result [36]) );
  dp_1 \pipeline/md/result_reg[37]  ( .ip(n8597), .ck(clk), .q(
        \pipeline/md/result [37]) );
  dp_1 \pipeline/md/result_reg[38]  ( .ip(n8596), .ck(clk), .q(
        \pipeline/md/result [38]) );
  dp_1 \pipeline/md/result_reg[39]  ( .ip(n8595), .ck(clk), .q(
        \pipeline/md/result [39]) );
  dp_1 \pipeline/md/result_reg[40]  ( .ip(n8594), .ck(clk), .q(
        \pipeline/md/result [40]) );
  dp_1 \pipeline/md/result_reg[41]  ( .ip(n8593), .ck(clk), .q(
        \pipeline/md/result [41]) );
  dp_1 \pipeline/md/result_reg[42]  ( .ip(n8592), .ck(clk), .q(
        \pipeline/md/result [42]) );
  dp_1 \pipeline/md/result_reg[43]  ( .ip(n8591), .ck(clk), .q(
        \pipeline/md/result [43]) );
  dp_1 \pipeline/md/result_reg[44]  ( .ip(n8590), .ck(clk), .q(
        \pipeline/md/result [44]) );
  dp_1 \pipeline/md/result_reg[45]  ( .ip(n8589), .ck(clk), .q(
        \pipeline/md/result [45]) );
  dp_1 \pipeline/md/result_reg[46]  ( .ip(n8588), .ck(clk), .q(
        \pipeline/md/result [46]) );
  dp_1 \pipeline/md/result_reg[47]  ( .ip(n8587), .ck(clk), .q(
        \pipeline/md/result [47]) );
  dp_1 \pipeline/md/result_reg[48]  ( .ip(n8586), .ck(clk), .q(
        \pipeline/md/result [48]) );
  dp_1 \pipeline/md/result_reg[49]  ( .ip(n8585), .ck(clk), .q(
        \pipeline/md/result [49]) );
  dp_1 \pipeline/md/result_reg[50]  ( .ip(n8584), .ck(clk), .q(
        \pipeline/md/result [50]) );
  dp_1 \pipeline/md/result_reg[51]  ( .ip(n8583), .ck(clk), .q(
        \pipeline/md/result [51]) );
  dp_1 \pipeline/md/result_reg[52]  ( .ip(n8582), .ck(clk), .q(
        \pipeline/md/result [52]) );
  dp_1 \pipeline/md/result_reg[53]  ( .ip(n8581), .ck(clk), .q(
        \pipeline/md/result [53]) );
  dp_1 \pipeline/md/result_reg[54]  ( .ip(n8580), .ck(clk), .q(
        \pipeline/md/result [54]) );
  dp_1 \pipeline/md/result_reg[55]  ( .ip(n8579), .ck(clk), .q(
        \pipeline/md/result [55]) );
  dp_1 \pipeline/md/result_reg[56]  ( .ip(n8578), .ck(clk), .q(
        \pipeline/md/result [56]) );
  dp_1 \pipeline/md/result_reg[57]  ( .ip(n8577), .ck(clk), .q(
        \pipeline/md/result [57]) );
  dp_1 \pipeline/md/result_reg[58]  ( .ip(n8576), .ck(clk), .q(
        \pipeline/md/result [58]) );
  dp_1 \pipeline/md/result_reg[59]  ( .ip(n8575), .ck(clk), .q(
        \pipeline/md/result [59]) );
  dp_1 \pipeline/md/result_reg[60]  ( .ip(n8574), .ck(clk), .q(
        \pipeline/md/result [60]) );
  dp_1 \pipeline/md/result_reg[61]  ( .ip(n8573), .ck(clk), .q(
        \pipeline/md/result [61]) );
  dp_1 \pipeline/md/result_reg[62]  ( .ip(n8572), .ck(clk), .q(
        \pipeline/md/result [62]) );
  dp_1 \pipeline/md/result_reg[63]  ( .ip(n8571), .ck(clk), .q(
        \pipeline/md/result [63]) );
  dp_1 \pipeline/md/a_reg[32]  ( .ip(n8570), .ck(clk), .q(\pipeline/md/a [32])
         );
  dp_1 \pipeline/md/a_reg[33]  ( .ip(n8569), .ck(clk), .q(\pipeline/md/a [33])
         );
  dp_1 \pipeline/md/a_reg[34]  ( .ip(n8568), .ck(clk), .q(\pipeline/md/a [34])
         );
  dp_1 \pipeline/md/a_reg[35]  ( .ip(n8567), .ck(clk), .q(\pipeline/md/a [35])
         );
  dp_1 \pipeline/md/a_reg[36]  ( .ip(n8566), .ck(clk), .q(\pipeline/md/a [36])
         );
  dp_1 \pipeline/md/a_reg[37]  ( .ip(n8565), .ck(clk), .q(\pipeline/md/a [37])
         );
  dp_1 \pipeline/md/a_reg[38]  ( .ip(n8564), .ck(clk), .q(\pipeline/md/a [38])
         );
  dp_1 \pipeline/md/a_reg[39]  ( .ip(n8563), .ck(clk), .q(\pipeline/md/a [39])
         );
  dp_1 \pipeline/md/a_reg[40]  ( .ip(n8562), .ck(clk), .q(\pipeline/md/a [40])
         );
  dp_1 \pipeline/md/a_reg[41]  ( .ip(n8561), .ck(clk), .q(\pipeline/md/a [41])
         );
  dp_1 \pipeline/md/a_reg[42]  ( .ip(n8560), .ck(clk), .q(\pipeline/md/a [42])
         );
  dp_1 \pipeline/md/a_reg[43]  ( .ip(n8559), .ck(clk), .q(\pipeline/md/a [43])
         );
  dp_1 \pipeline/md/a_reg[44]  ( .ip(n8558), .ck(clk), .q(\pipeline/md/a [44])
         );
  dp_1 \pipeline/md/a_reg[45]  ( .ip(n8557), .ck(clk), .q(\pipeline/md/a [45])
         );
  dp_1 \pipeline/md/a_reg[46]  ( .ip(n8556), .ck(clk), .q(\pipeline/md/a [46])
         );
  dp_1 \pipeline/md/a_reg[47]  ( .ip(n8555), .ck(clk), .q(\pipeline/md/a [47])
         );
  dp_1 \pipeline/md/a_reg[48]  ( .ip(n8554), .ck(clk), .q(\pipeline/md/a [48])
         );
  dp_1 \pipeline/md/a_reg[49]  ( .ip(n8553), .ck(clk), .q(\pipeline/md/a [49])
         );
  dp_1 \pipeline/md/a_reg[50]  ( .ip(n8552), .ck(clk), .q(\pipeline/md/a [50])
         );
  dp_1 \pipeline/md/a_reg[51]  ( .ip(n8551), .ck(clk), .q(\pipeline/md/a [51])
         );
  dp_1 \pipeline/md/a_reg[52]  ( .ip(n8550), .ck(clk), .q(\pipeline/md/a [52])
         );
  dp_1 \pipeline/md/a_reg[53]  ( .ip(n8549), .ck(clk), .q(\pipeline/md/a [53])
         );
  dp_1 \pipeline/md/a_reg[54]  ( .ip(n8548), .ck(clk), .q(\pipeline/md/a [54])
         );
  dp_1 \pipeline/md/a_reg[55]  ( .ip(n8547), .ck(clk), .q(\pipeline/md/a [55])
         );
  dp_1 \pipeline/md/a_reg[56]  ( .ip(n8546), .ck(clk), .q(\pipeline/md/a [56])
         );
  dp_1 \pipeline/md/a_reg[57]  ( .ip(n8545), .ck(clk), .q(\pipeline/md/a [57])
         );
  dp_1 \pipeline/md/a_reg[58]  ( .ip(n8544), .ck(clk), .q(\pipeline/md/a [58])
         );
  dp_1 \pipeline/md/a_reg[59]  ( .ip(n8543), .ck(clk), .q(\pipeline/md/a [59])
         );
  dp_1 \pipeline/md/a_reg[60]  ( .ip(n8542), .ck(clk), .q(\pipeline/md/a [60])
         );
  dp_1 \pipeline/md/a_reg[61]  ( .ip(n8541), .ck(clk), .q(\pipeline/md/a [61])
         );
  dp_1 \pipeline/md/a_reg[62]  ( .ip(n8540), .ck(clk), .q(\pipeline/md/a [62])
         );
  dp_1 \pipeline/md/counter_reg[0]  ( .ip(n8538), .ck(clk), .q(
        \pipeline/md/counter [0]) );
  dp_1 \pipeline/md/counter_reg[1]  ( .ip(n8537), .ck(clk), .q(
        \pipeline/md/counter [1]) );
  dp_1 \pipeline/md/counter_reg[2]  ( .ip(n8536), .ck(clk), .q(
        \pipeline/md/counter [2]) );
  dp_1 \pipeline/md/counter_reg[3]  ( .ip(n8535), .ck(clk), .q(
        \pipeline/md/counter [3]) );
  dp_1 \pipeline/md/counter_reg[4]  ( .ip(n8534), .ck(clk), .q(
        \pipeline/md/counter [4]) );
  dp_1 \pipeline/inst_DX_reg[2]  ( .ip(n8533), .ck(clk), .q(
        \pipeline/inst_DX [2]) );
  dp_1 \pipeline/inst_DX_reg[3]  ( .ip(n8532), .ck(clk), .q(
        \pipeline/inst_DX [3]) );
  dp_1 \pipeline/inst_DX_reg[5]  ( .ip(n8531), .ck(clk), .q(
        \pipeline/inst_DX [5]) );
  dp_1 \pipeline/inst_DX_reg[6]  ( .ip(n8530), .ck(clk), .q(
        \pipeline/inst_DX [6]) );
  dp_1 \pipeline/inst_DX_reg[7]  ( .ip(n8529), .ck(clk), .q(
        \pipeline/inst_DX [7]) );
  dp_1 \pipeline/inst_DX_reg[8]  ( .ip(n8528), .ck(clk), .q(
        \pipeline/inst_DX [8]) );
  dp_1 \pipeline/inst_DX_reg[9]  ( .ip(n8527), .ck(clk), .q(
        \pipeline/inst_DX [9]) );
  dp_1 \pipeline/inst_DX_reg[10]  ( .ip(n8526), .ck(clk), .q(
        \pipeline/inst_DX [10]) );
  dp_1 \pipeline/inst_DX_reg[11]  ( .ip(n8525), .ck(clk), .q(
        \pipeline/inst_DX [11]) );
  dp_1 \pipeline/md/a_reg[31]  ( .ip(n8521), .ck(clk), .q(\pipeline/md/a [31])
         );
  dp_1 \pipeline/inst_DX_reg[15]  ( .ip(n8520), .ck(clk), .q(
        \pipeline/inst_DX [15]) );
  dp_1 \pipeline/inst_DX_reg[16]  ( .ip(n8519), .ck(clk), .q(
        \pipeline/inst_DX [16]) );
  dp_1 \pipeline/inst_DX_reg[18]  ( .ip(n8517), .ck(clk), .q(
        \pipeline/inst_DX [18]) );
  dp_1 \pipeline/inst_DX_reg[19]  ( .ip(n8516), .ck(clk), .q(
        \pipeline/inst_DX [19]) );
  dp_1 \pipeline/inst_DX_reg[20]  ( .ip(n8515), .ck(clk), .q(
        \pipeline/inst_DX [20]) );
  dp_1 \pipeline/inst_DX_reg[21]  ( .ip(n8514), .ck(clk), .q(
        \pipeline/inst_DX [21]) );
  dp_1 \pipeline/inst_DX_reg[23]  ( .ip(n8512), .ck(clk), .q(
        \pipeline/inst_DX [23]) );
  dp_1 \pipeline/inst_DX_reg[24]  ( .ip(n8511), .ck(clk), .q(
        \pipeline/inst_DX [24]) );
  dp_1 \pipeline/inst_DX_reg[25]  ( .ip(n8510), .ck(clk), .q(
        \pipeline/inst_DX [25]) );
  dp_1 \pipeline/inst_DX_reg[28]  ( .ip(n8507), .ck(clk), .q(
        \pipeline/inst_DX [28]) );
  dp_1 \pipeline/inst_DX_reg[29]  ( .ip(n8506), .ck(clk), .q(
        \pipeline/inst_DX [29]) );
  dp_1 \pipeline/inst_DX_reg[31]  ( .ip(n8504), .ck(clk), .q(
        \pipeline/imm[31] ) );
  dp_1 \pipeline/inst_DX_reg[0]  ( .ip(n8503), .ck(clk), .q(
        \pipeline/inst_DX [0]) );
  dp_1 \pipeline/inst_DX_reg[1]  ( .ip(n8502), .ck(clk), .q(
        \pipeline/inst_DX [1]) );
  dp_1 \pipeline/inst_DX_reg[4]  ( .ip(n8501), .ck(clk), .q(
        \pipeline/inst_DX [4]) );
  dp_1 \pipeline/ctrl/had_ex_DX_reg  ( .ip(n8500), .ck(clk), .q(
        \pipeline/ctrl/had_ex_DX ) );
  dp_1 \pipeline/ctrl/had_ex_WB_reg  ( .ip(n8499), .ck(clk), .q(
        \pipeline/ctrl/had_ex_WB ) );
  dp_1 \pipeline/ctrl/store_in_WB_reg  ( .ip(n8498), .ck(clk), .q(
        \pipeline/ctrl/store_in_WB ) );
  dp_1 \pipeline/ctrl/dmem_en_WB_reg  ( .ip(n8497), .ck(clk), .q(
        \pipeline/ctrl/dmem_en_WB ) );
  dp_1 \pipeline/md/b_reg[62]  ( .ip(n8496), .ck(clk), .q(\pipeline/md/b [62])
         );
  dp_1 \pipeline/ctrl/wr_reg_unkilled_WB_reg  ( .ip(n8495), .ck(clk), .q(
        \pipeline/ctrl/wr_reg_unkilled_WB ) );
  dp_1 \pipeline/ctrl/wfi_unkilled_WB_reg  ( .ip(n8494), .ck(clk), .q(
        \pipeline/ctrl/wfi_unkilled_WB ) );
  dp_1 \pipeline/ctrl/uses_md_WB_reg  ( .ip(n8493), .ck(clk), .q(
        \pipeline/ctrl/uses_md_WB ) );
  dp_1 \pipeline/ctrl/prev_killed_DX_reg  ( .ip(n8492), .ck(clk), .q(
        \pipeline/ctrl/prev_killed_DX ) );
  dp_1 \pipeline/ctrl/prev_killed_WB_reg  ( .ip(n8491), .ck(clk), .q(
        \pipeline/ctrl/prev_killed_WB ) );
  dp_1 \pipeline/PC_IF_reg[0]  ( .ip(n8490), .ck(clk), .q(\pipeline/PC_IF [0])
         );
  dp_1 \pipeline/PC_DX_reg[0]  ( .ip(n8489), .ck(clk), .q(\pipeline/PC_DX [0])
         );
  dp_1 \pipeline/PC_IF_reg[1]  ( .ip(n8488), .ck(clk), .q(\pipeline/PC_IF [1])
         );
  dp_1 \pipeline/PC_DX_reg[1]  ( .ip(n8487), .ck(clk), .q(\pipeline/PC_DX [1])
         );
  dp_1 \pipeline/PC_IF_reg[2]  ( .ip(n8486), .ck(clk), .q(\pipeline/PC_IF [2])
         );
  dp_1 \pipeline/PC_DX_reg[2]  ( .ip(n8485), .ck(clk), .q(\pipeline/PC_DX [2])
         );
  dp_1 \pipeline/PC_IF_reg[3]  ( .ip(n8484), .ck(clk), .q(\pipeline/PC_IF [3])
         );
  dp_1 \pipeline/PC_DX_reg[3]  ( .ip(n8483), .ck(clk), .q(\pipeline/PC_DX [3])
         );
  dp_1 \pipeline/PC_IF_reg[4]  ( .ip(n8482), .ck(clk), .q(\pipeline/PC_IF [4])
         );
  dp_1 \pipeline/PC_DX_reg[4]  ( .ip(n8481), .ck(clk), .q(\pipeline/PC_DX [4])
         );
  dp_1 \pipeline/PC_IF_reg[5]  ( .ip(n8480), .ck(clk), .q(\pipeline/PC_IF [5])
         );
  dp_1 \pipeline/PC_DX_reg[5]  ( .ip(n8479), .ck(clk), .q(\pipeline/PC_DX [5])
         );
  dp_1 \pipeline/PC_IF_reg[6]  ( .ip(n8478), .ck(clk), .q(\pipeline/PC_IF [6])
         );
  dp_1 \pipeline/PC_DX_reg[6]  ( .ip(n8477), .ck(clk), .q(\pipeline/PC_DX [6])
         );
  dp_1 \pipeline/PC_IF_reg[7]  ( .ip(n8476), .ck(clk), .q(\pipeline/PC_IF [7])
         );
  dp_1 \pipeline/PC_DX_reg[7]  ( .ip(n8475), .ck(clk), .q(\pipeline/PC_DX [7])
         );
  dp_1 \pipeline/PC_IF_reg[8]  ( .ip(n8474), .ck(clk), .q(\pipeline/PC_IF [8])
         );
  dp_1 \pipeline/PC_DX_reg[8]  ( .ip(n8473), .ck(clk), .q(\pipeline/PC_DX [8])
         );
  dp_1 \pipeline/PC_IF_reg[9]  ( .ip(n8472), .ck(clk), .q(\pipeline/PC_IF [9])
         );
  dp_1 \pipeline/PC_DX_reg[9]  ( .ip(n8471), .ck(clk), .q(\pipeline/PC_DX [9])
         );
  dp_1 \pipeline/PC_IF_reg[10]  ( .ip(n8470), .ck(clk), .q(
        \pipeline/PC_IF [10]) );
  dp_1 \pipeline/PC_DX_reg[10]  ( .ip(n8469), .ck(clk), .q(
        \pipeline/PC_DX [10]) );
  dp_1 \pipeline/PC_IF_reg[11]  ( .ip(n8468), .ck(clk), .q(
        \pipeline/PC_IF [11]) );
  dp_1 \pipeline/PC_DX_reg[11]  ( .ip(n8467), .ck(clk), .q(
        \pipeline/PC_DX [11]) );
  dp_1 \pipeline/PC_IF_reg[12]  ( .ip(n8466), .ck(clk), .q(
        \pipeline/PC_IF [12]) );
  dp_1 \pipeline/PC_DX_reg[12]  ( .ip(n8465), .ck(clk), .q(
        \pipeline/PC_DX [12]) );
  dp_1 \pipeline/PC_IF_reg[13]  ( .ip(n8464), .ck(clk), .q(
        \pipeline/PC_IF [13]) );
  dp_1 \pipeline/PC_DX_reg[13]  ( .ip(n8463), .ck(clk), .q(
        \pipeline/PC_DX [13]) );
  dp_1 \pipeline/PC_IF_reg[14]  ( .ip(n8462), .ck(clk), .q(
        \pipeline/PC_IF [14]) );
  dp_1 \pipeline/PC_DX_reg[14]  ( .ip(n8461), .ck(clk), .q(
        \pipeline/PC_DX [14]) );
  dp_1 \pipeline/PC_IF_reg[15]  ( .ip(n8460), .ck(clk), .q(
        \pipeline/PC_IF [15]) );
  dp_1 \pipeline/PC_DX_reg[15]  ( .ip(n8459), .ck(clk), .q(
        \pipeline/PC_DX [15]) );
  dp_1 \pipeline/PC_IF_reg[16]  ( .ip(n8458), .ck(clk), .q(
        \pipeline/PC_IF [16]) );
  dp_1 \pipeline/PC_DX_reg[16]  ( .ip(n8457), .ck(clk), .q(
        \pipeline/PC_DX [16]) );
  dp_1 \pipeline/PC_IF_reg[17]  ( .ip(n8456), .ck(clk), .q(
        \pipeline/PC_IF [17]) );
  dp_1 \pipeline/PC_DX_reg[17]  ( .ip(n8455), .ck(clk), .q(
        \pipeline/PC_DX [17]) );
  dp_1 \pipeline/PC_IF_reg[18]  ( .ip(n8454), .ck(clk), .q(
        \pipeline/PC_IF [18]) );
  dp_1 \pipeline/PC_DX_reg[18]  ( .ip(n8453), .ck(clk), .q(
        \pipeline/PC_DX [18]) );
  dp_1 \pipeline/PC_IF_reg[19]  ( .ip(n8452), .ck(clk), .q(
        \pipeline/PC_IF [19]) );
  dp_1 \pipeline/PC_DX_reg[19]  ( .ip(n8451), .ck(clk), .q(
        \pipeline/PC_DX [19]) );
  dp_1 \pipeline/PC_IF_reg[20]  ( .ip(n8450), .ck(clk), .q(
        \pipeline/PC_IF [20]) );
  dp_1 \pipeline/PC_DX_reg[20]  ( .ip(n8449), .ck(clk), .q(
        \pipeline/PC_DX [20]) );
  dp_1 \pipeline/PC_IF_reg[21]  ( .ip(n8448), .ck(clk), .q(
        \pipeline/PC_IF [21]) );
  dp_1 \pipeline/PC_DX_reg[21]  ( .ip(n8447), .ck(clk), .q(
        \pipeline/PC_DX [21]) );
  dp_1 \pipeline/PC_IF_reg[22]  ( .ip(n8446), .ck(clk), .q(
        \pipeline/PC_IF [22]) );
  dp_1 \pipeline/PC_DX_reg[22]  ( .ip(n8445), .ck(clk), .q(
        \pipeline/PC_DX [22]) );
  dp_1 \pipeline/PC_IF_reg[23]  ( .ip(n8444), .ck(clk), .q(
        \pipeline/PC_IF [23]) );
  dp_1 \pipeline/PC_DX_reg[23]  ( .ip(n8443), .ck(clk), .q(
        \pipeline/PC_DX [23]) );
  dp_1 \pipeline/PC_IF_reg[24]  ( .ip(n8442), .ck(clk), .q(
        \pipeline/PC_IF [24]) );
  dp_1 \pipeline/PC_DX_reg[24]  ( .ip(n8441), .ck(clk), .q(
        \pipeline/PC_DX [24]) );
  dp_1 \pipeline/PC_IF_reg[25]  ( .ip(n8440), .ck(clk), .q(
        \pipeline/PC_IF [25]) );
  dp_1 \pipeline/PC_DX_reg[25]  ( .ip(n8439), .ck(clk), .q(
        \pipeline/PC_DX [25]) );
  dp_1 \pipeline/PC_IF_reg[26]  ( .ip(n8438), .ck(clk), .q(
        \pipeline/PC_IF [26]) );
  dp_1 \pipeline/PC_DX_reg[26]  ( .ip(n8437), .ck(clk), .q(
        \pipeline/PC_DX [26]) );
  dp_1 \pipeline/PC_IF_reg[27]  ( .ip(n8436), .ck(clk), .q(
        \pipeline/PC_IF [27]) );
  dp_1 \pipeline/PC_DX_reg[27]  ( .ip(n8435), .ck(clk), .q(
        \pipeline/PC_DX [27]) );
  dp_1 \pipeline/PC_IF_reg[28]  ( .ip(n8434), .ck(clk), .q(
        \pipeline/PC_IF [28]) );
  dp_1 \pipeline/PC_DX_reg[28]  ( .ip(n8433), .ck(clk), .q(
        \pipeline/PC_DX [28]) );
  dp_1 \pipeline/PC_IF_reg[29]  ( .ip(n8432), .ck(clk), .q(
        \pipeline/PC_IF [29]) );
  dp_1 \pipeline/PC_DX_reg[29]  ( .ip(n8431), .ck(clk), .q(
        \pipeline/PC_DX [29]) );
  dp_1 \pipeline/PC_IF_reg[30]  ( .ip(n8430), .ck(clk), .q(
        \pipeline/PC_IF [30]) );
  dp_1 \pipeline/PC_DX_reg[30]  ( .ip(n8429), .ck(clk), .q(
        \pipeline/PC_DX [30]) );
  dp_1 \pipeline/PC_IF_reg[31]  ( .ip(n8428), .ck(clk), .q(
        \pipeline/PC_IF [31]) );
  dp_1 \pipeline/PC_DX_reg[31]  ( .ip(n8427), .ck(clk), .q(
        \pipeline/PC_DX [31]) );
  dp_1 \pipeline/md/a_reg[0]  ( .ip(n8426), .ck(clk), .q(\pipeline/md/a [0])
         );
  dp_1 \pipeline/md/a_reg[16]  ( .ip(n8425), .ck(clk), .q(\pipeline/md/a [16])
         );
  dp_1 \pipeline/md/a_reg[24]  ( .ip(n8424), .ck(clk), .q(\pipeline/md/a [24])
         );
  dp_1 \pipeline/md/a_reg[28]  ( .ip(n8423), .ck(clk), .q(\pipeline/md/a [28])
         );
  dp_1 \pipeline/md/b_reg[61]  ( .ip(n8422), .ck(clk), .q(\pipeline/md/b [61])
         );
  dp_1 \pipeline/md/a_reg[30]  ( .ip(n8421), .ck(clk), .q(\pipeline/md/a [30])
         );
  dp_1 \pipeline/md/a_reg[11]  ( .ip(n8420), .ck(clk), .q(\pipeline/md/a [11])
         );
  dp_1 \pipeline/md/a_reg[27]  ( .ip(n8419), .ck(clk), .q(\pipeline/md/a [27])
         );
  dp_1 \pipeline/md/b_reg[60]  ( .ip(n8418), .ck(clk), .q(\pipeline/md/b [60])
         );
  dp_1 \pipeline/md/b_reg[59]  ( .ip(n8417), .ck(clk), .q(\pipeline/md/b [59])
         );
  dp_1 \pipeline/md/b_reg[58]  ( .ip(n8416), .ck(clk), .q(\pipeline/md/b [58])
         );
  dp_1 \pipeline/md/a_reg[29]  ( .ip(n8415), .ck(clk), .q(\pipeline/md/a [29])
         );
  dp_1 \pipeline/md/a_reg[10]  ( .ip(n8414), .ck(clk), .q(\pipeline/md/a [10])
         );
  dp_1 \pipeline/md/b_reg[57]  ( .ip(n8413), .ck(clk), .q(\pipeline/md/b [57])
         );
  dp_1 \pipeline/md/a_reg[26]  ( .ip(n8412), .ck(clk), .q(\pipeline/md/a [26])
         );
  dp_1 \pipeline/md/a_reg[12]  ( .ip(n8411), .ck(clk), .q(\pipeline/md/a [12])
         );
  dp_1 \pipeline/md/a_reg[20]  ( .ip(n8410), .ck(clk), .q(\pipeline/md/a [20])
         );
  dp_1 \pipeline/md/a_reg[22]  ( .ip(n8409), .ck(clk), .q(\pipeline/md/a [22])
         );
  dp_1 \pipeline/md/a_reg[23]  ( .ip(n8408), .ck(clk), .q(\pipeline/md/a [23])
         );
  dp_1 \pipeline/md/a_reg[8]  ( .ip(n8407), .ck(clk), .q(\pipeline/md/a [8])
         );
  dp_1 \pipeline/md/a_reg[13]  ( .ip(n8406), .ck(clk), .q(\pipeline/md/a [13])
         );
  dp_1 \pipeline/md/a_reg[17]  ( .ip(n8405), .ck(clk), .q(\pipeline/md/a [17])
         );
  dp_1 \pipeline/md/a_reg[21]  ( .ip(n8404), .ck(clk), .q(\pipeline/md/a [21])
         );
  dp_1 \pipeline/md/b_reg[56]  ( .ip(n8403), .ck(clk), .q(\pipeline/md/b [56])
         );
  dp_1 \pipeline/md/b_reg[55]  ( .ip(n8402), .ck(clk), .q(\pipeline/md/b [55])
         );
  dp_1 \pipeline/md/b_reg[54]  ( .ip(n22861), .ck(clk), .q(\pipeline/md/b [54]) );
  dp_1 \pipeline/md/b_reg[53]  ( .ip(n8400), .ck(clk), .q(\pipeline/md/b [53])
         );
  dp_1 \pipeline/md/b_reg[52]  ( .ip(n22860), .ck(clk), .q(\pipeline/md/b [52]) );
  dp_1 \pipeline/md/b_reg[51]  ( .ip(n8398), .ck(clk), .q(\pipeline/md/b [51])
         );
  dp_1 \pipeline/md/a_reg[25]  ( .ip(n8397), .ck(clk), .q(\pipeline/md/a [25])
         );
  dp_1 \pipeline/md/a_reg[18]  ( .ip(n8396), .ck(clk), .q(\pipeline/md/a [18])
         );
  dp_1 \pipeline/md/b_reg[50]  ( .ip(n8395), .ck(clk), .q(\pipeline/md/b [50])
         );
  dp_1 \pipeline/md/b_reg[49]  ( .ip(n8394), .ck(clk), .q(\pipeline/md/b [49])
         );
  dp_1 \pipeline/md/b_reg[48]  ( .ip(n8393), .ck(clk), .q(\pipeline/md/b [48])
         );
  dp_1 \pipeline/md/b_reg[47]  ( .ip(n8392), .ck(clk), .q(\pipeline/md/b [47])
         );
  dp_1 \pipeline/md/a_reg[19]  ( .ip(n8391), .ck(clk), .q(\pipeline/md/a [19])
         );
  dp_1 \pipeline/md/a_reg[4]  ( .ip(n8390), .ck(clk), .q(\pipeline/md/a [4])
         );
  dp_1 \pipeline/md/a_reg[14]  ( .ip(n8389), .ck(clk), .q(\pipeline/md/a [14])
         );
  dp_1 \pipeline/md/b_reg[46]  ( .ip(n22859), .ck(clk), .q(\pipeline/md/b [46]) );
  dp_1 \pipeline/md/b_reg[45]  ( .ip(n8387), .ck(clk), .q(\pipeline/md/b [45])
         );
  dp_1 \pipeline/md/b_reg[44]  ( .ip(n8386), .ck(clk), .q(\pipeline/md/b [44])
         );
  dp_1 \pipeline/md/b_reg[43]  ( .ip(n8385), .ck(clk), .q(\pipeline/md/b [43])
         );
  dp_1 \pipeline/md/b_reg[42]  ( .ip(n8384), .ck(clk), .q(\pipeline/md/b [42])
         );
  dp_1 \pipeline/md/b_reg[41]  ( .ip(n22862), .ck(clk), .q(\pipeline/md/b [41]) );
  dp_1 \pipeline/md/a_reg[15]  ( .ip(n8382), .ck(clk), .q(\pipeline/md/a [15])
         );
  dp_1 \pipeline/md/a_reg[2]  ( .ip(n22855), .ck(clk), .q(\pipeline/md/a [2])
         );
  dp_1 \pipeline/md/a_reg[3]  ( .ip(n8380), .ck(clk), .q(\pipeline/md/a [3])
         );
  dp_1 \pipeline/md/a_reg[1]  ( .ip(n22854), .ck(clk), .q(\pipeline/md/a [1])
         );
  dp_1 \pipeline/md/a_reg[5]  ( .ip(n8378), .ck(clk), .q(\pipeline/md/a [5])
         );
  dp_1 \pipeline/md/b_reg[40]  ( .ip(n8377), .ck(clk), .q(\pipeline/md/b [40])
         );
  dp_1 \pipeline/md/b_reg[39]  ( .ip(n8376), .ck(clk), .q(\pipeline/md/b [39])
         );
  dp_1 \pipeline/md/a_reg[9]  ( .ip(n8375), .ck(clk), .q(\pipeline/md/a [9])
         );
  dp_1 \pipeline/md/b_reg[38]  ( .ip(n8374), .ck(clk), .q(\pipeline/md/b [38])
         );
  dp_1 \pipeline/md/a_reg[7]  ( .ip(n8373), .ck(clk), .q(\pipeline/md/a [7])
         );
  dp_1 \pipeline/md/b_reg[37]  ( .ip(n8372), .ck(clk), .q(\pipeline/md/b [37])
         );
  dp_1 \pipeline/md/b_reg[36]  ( .ip(n8371), .ck(clk), .q(\pipeline/md/b [36])
         );
  dp_1 \pipeline/md/b_reg[35]  ( .ip(n22850), .ck(clk), .q(\pipeline/md/b [35]) );
  dp_1 \pipeline/md/b_reg[34]  ( .ip(n8369), .ck(clk), .q(\pipeline/md/b [34])
         );
  dp_1 \pipeline/md/b_reg[33]  ( .ip(n8368), .ck(clk), .q(\pipeline/md/b [33])
         );
  dp_1 \pipeline/md/b_reg[32]  ( .ip(n8367), .ck(clk), .q(\pipeline/md/b [32])
         );
  dp_1 \pipeline/md/a_reg[6]  ( .ip(n8366), .ck(clk), .q(\pipeline/md/a [6])
         );
  dp_1 \pipeline/md/b_reg[31]  ( .ip(n8365), .ck(clk), .q(\pipeline/md/b [31])
         );
  dp_1 \pipeline/md/b_reg[30]  ( .ip(n8364), .ck(clk), .q(\pipeline/md/b [30])
         );
  dp_1 \pipeline/md/b_reg[29]  ( .ip(n8363), .ck(clk), .q(\pipeline/md/b [29])
         );
  dp_1 \pipeline/md/b_reg[28]  ( .ip(n8362), .ck(clk), .q(\pipeline/md/b [28])
         );
  dp_1 \pipeline/md/b_reg[27]  ( .ip(n8361), .ck(clk), .q(\pipeline/md/b [27])
         );
  dp_1 \pipeline/md/b_reg[26]  ( .ip(n8360), .ck(clk), .q(\pipeline/md/b [26])
         );
  dp_1 \pipeline/md/b_reg[25]  ( .ip(n8359), .ck(clk), .q(\pipeline/md/b [25])
         );
  dp_1 \pipeline/md/b_reg[24]  ( .ip(n8358), .ck(clk), .q(\pipeline/md/b [24])
         );
  dp_1 \pipeline/md/b_reg[23]  ( .ip(n8357), .ck(clk), .q(\pipeline/md/b [23])
         );
  dp_1 \pipeline/md/b_reg[22]  ( .ip(n8356), .ck(clk), .q(\pipeline/md/b [22])
         );
  dp_1 \pipeline/md/b_reg[21]  ( .ip(n8355), .ck(clk), .q(\pipeline/md/b [21])
         );
  dp_1 \pipeline/md/b_reg[20]  ( .ip(n8354), .ck(clk), .q(\pipeline/md/b [20])
         );
  dp_1 \pipeline/md/b_reg[19]  ( .ip(n8353), .ck(clk), .q(\pipeline/md/b [19])
         );
  dp_1 \pipeline/md/b_reg[18]  ( .ip(n8352), .ck(clk), .q(\pipeline/md/b [18])
         );
  dp_1 \pipeline/md/b_reg[17]  ( .ip(n8351), .ck(clk), .q(\pipeline/md/b [17])
         );
  dp_1 \pipeline/md/b_reg[16]  ( .ip(n8350), .ck(clk), .q(\pipeline/md/b [16])
         );
  dp_1 \pipeline/md/b_reg[15]  ( .ip(n8349), .ck(clk), .q(\pipeline/md/b [15])
         );
  dp_1 \pipeline/md/b_reg[14]  ( .ip(n8348), .ck(clk), .q(\pipeline/md/b [14])
         );
  dp_1 \pipeline/md/b_reg[13]  ( .ip(n8347), .ck(clk), .q(\pipeline/md/b [13])
         );
  dp_1 \pipeline/md/b_reg[12]  ( .ip(n8346), .ck(clk), .q(\pipeline/md/b [12])
         );
  dp_1 \pipeline/md/b_reg[11]  ( .ip(n8345), .ck(clk), .q(\pipeline/md/b [11])
         );
  dp_1 \pipeline/md/b_reg[10]  ( .ip(n8344), .ck(clk), .q(\pipeline/md/b [10])
         );
  dp_1 \pipeline/md/b_reg[9]  ( .ip(n8343), .ck(clk), .q(\pipeline/md/b [9])
         );
  dp_1 \pipeline/md/b_reg[8]  ( .ip(n8342), .ck(clk), .q(\pipeline/md/b [8])
         );
  dp_1 \pipeline/md/b_reg[7]  ( .ip(n8341), .ck(clk), .q(\pipeline/md/b [7])
         );
  dp_1 \pipeline/md/b_reg[6]  ( .ip(n8340), .ck(clk), .q(\pipeline/md/b [6])
         );
  dp_1 \pipeline/md/b_reg[5]  ( .ip(n8339), .ck(clk), .q(\pipeline/md/b [5])
         );
  dp_1 \pipeline/md/b_reg[4]  ( .ip(n8338), .ck(clk), .q(\pipeline/md/b [4])
         );
  dp_1 \pipeline/md/b_reg[3]  ( .ip(n8337), .ck(clk), .q(\pipeline/md/b [3])
         );
  dp_1 \pipeline/md/b_reg[2]  ( .ip(n8336), .ck(clk), .q(\pipeline/md/b [2])
         );
  dp_1 \pipeline/md/b_reg[1]  ( .ip(n8335), .ck(clk), .q(\pipeline/md/b [1])
         );
  dp_1 \pipeline/md/b_reg[0]  ( .ip(n8334), .ck(clk), .q(\pipeline/md/b [0])
         );
  dp_1 \pipeline/md/state_reg[0]  ( .ip(n17756), .ck(clk), .q(
        \pipeline/md/state [0]) );
  dp_1 \pipeline/md/state_reg[1]  ( .ip(\pipeline/md/N162 ), .ck(clk), .q(
        \pipeline/md/state [1]) );
  dp_1 \pipeline/csr/htif_state_reg  ( .ip(n10139), .ck(clk), .q(
        htif_pcr_resp_valid) );
  dp_1 \pipeline/csr/to_host_reg[0]  ( .ip(n8772), .ck(clk), .q(
        \pipeline/csr/to_host [0]) );
  dp_1 \pipeline/csr/to_host_reg[1]  ( .ip(n8771), .ck(clk), .q(
        \pipeline/csr/to_host [1]) );
  dp_1 \pipeline/csr/to_host_reg[2]  ( .ip(n8770), .ck(clk), .q(
        \pipeline/csr/to_host [2]) );
  dp_1 \pipeline/csr/to_host_reg[3]  ( .ip(n8769), .ck(clk), .q(
        \pipeline/csr/to_host [3]) );
  dp_1 \pipeline/csr/to_host_reg[4]  ( .ip(n8768), .ck(clk), .q(
        \pipeline/csr/to_host [4]) );
  dp_1 \pipeline/csr/to_host_reg[5]  ( .ip(n8767), .ck(clk), .q(
        \pipeline/csr/to_host [5]) );
  dp_1 \pipeline/csr/to_host_reg[6]  ( .ip(n8766), .ck(clk), .q(
        \pipeline/csr/to_host [6]) );
  dp_1 \pipeline/csr/to_host_reg[7]  ( .ip(n8765), .ck(clk), .q(
        \pipeline/csr/to_host [7]) );
  dp_1 \pipeline/csr/to_host_reg[8]  ( .ip(n8764), .ck(clk), .q(
        \pipeline/csr/to_host [8]) );
  dp_1 \pipeline/csr/to_host_reg[9]  ( .ip(n8763), .ck(clk), .q(
        \pipeline/csr/to_host [9]) );
  dp_1 \pipeline/csr/to_host_reg[10]  ( .ip(n8762), .ck(clk), .q(
        \pipeline/csr/to_host [10]) );
  dp_1 \pipeline/csr/to_host_reg[11]  ( .ip(n8761), .ck(clk), .q(
        \pipeline/csr/to_host [11]) );
  dp_1 \pipeline/csr/to_host_reg[12]  ( .ip(n8760), .ck(clk), .q(
        \pipeline/csr/to_host [12]) );
  dp_1 \pipeline/csr/to_host_reg[13]  ( .ip(n8759), .ck(clk), .q(
        \pipeline/csr/to_host [13]) );
  dp_1 \pipeline/csr/to_host_reg[14]  ( .ip(n8758), .ck(clk), .q(
        \pipeline/csr/to_host [14]) );
  dp_1 \pipeline/csr/to_host_reg[15]  ( .ip(n8757), .ck(clk), .q(
        \pipeline/csr/to_host [15]) );
  dp_1 \pipeline/csr/to_host_reg[16]  ( .ip(n8756), .ck(clk), .q(
        \pipeline/csr/to_host [16]) );
  dp_1 \pipeline/csr/to_host_reg[17]  ( .ip(n8755), .ck(clk), .q(
        \pipeline/csr/to_host [17]) );
  dp_1 \pipeline/csr/to_host_reg[18]  ( .ip(n8754), .ck(clk), .q(
        \pipeline/csr/to_host [18]) );
  dp_1 \pipeline/csr/to_host_reg[19]  ( .ip(n8753), .ck(clk), .q(
        \pipeline/csr/to_host [19]) );
  dp_1 \pipeline/csr/to_host_reg[20]  ( .ip(n8752), .ck(clk), .q(
        \pipeline/csr/to_host [20]) );
  dp_1 \pipeline/csr/to_host_reg[21]  ( .ip(n8751), .ck(clk), .q(
        \pipeline/csr/to_host [21]) );
  dp_1 \pipeline/csr/to_host_reg[22]  ( .ip(n8750), .ck(clk), .q(
        \pipeline/csr/to_host [22]) );
  dp_1 \pipeline/csr/to_host_reg[23]  ( .ip(n8749), .ck(clk), .q(
        \pipeline/csr/to_host [23]) );
  dp_1 \pipeline/csr/to_host_reg[24]  ( .ip(n8748), .ck(clk), .q(
        \pipeline/csr/to_host [24]) );
  dp_1 \pipeline/csr/to_host_reg[25]  ( .ip(n8747), .ck(clk), .q(
        \pipeline/csr/to_host [25]) );
  dp_1 \pipeline/csr/to_host_reg[26]  ( .ip(n8746), .ck(clk), .q(
        \pipeline/csr/to_host [26]) );
  dp_1 \pipeline/csr/to_host_reg[27]  ( .ip(n8745), .ck(clk), .q(
        \pipeline/csr/to_host [27]) );
  dp_1 \pipeline/csr/to_host_reg[28]  ( .ip(n8744), .ck(clk), .q(
        \pipeline/csr/to_host [28]) );
  dp_1 \pipeline/csr/to_host_reg[29]  ( .ip(n8743), .ck(clk), .q(
        \pipeline/csr/to_host [29]) );
  dp_1 \pipeline/csr/to_host_reg[30]  ( .ip(n8742), .ck(clk), .q(
        \pipeline/csr/to_host [30]) );
  dp_1 \pipeline/csr/to_host_reg[31]  ( .ip(n8741), .ck(clk), .q(
        \pipeline/csr/to_host [31]) );
  dp_1 \pipeline/csr_rdata_WB_reg[31]  ( .ip(n10072), .ck(clk), .q(
        \pipeline/csr_rdata_WB [31]) );
  dp_1 \pipeline/csr/msip_reg  ( .ip(n10074), .ck(clk), .q(
        \pipeline/csr/mip_3 ) );
  dp_1 \pipeline/csr/mtip_reg  ( .ip(n10073), .ck(clk), .q(
        \pipeline/csr/mip[7] ) );
  dp_1 \pipeline/ctrl/reg_to_wr_WB_reg[4]  ( .ip(n10071), .ck(clk), .q(
        \pipeline/reg_to_wr_WB [4]) );
  dp_1 \pipeline/ctrl/reg_to_wr_WB_reg[0]  ( .ip(n10070), .ck(clk), .q(
        \pipeline/reg_to_wr_WB [0]) );
  dp_1 \pipeline/ctrl/reg_to_wr_WB_reg[1]  ( .ip(n10069), .ck(clk), .q(
        \pipeline/reg_to_wr_WB [1]) );
  dp_1 \pipeline/ctrl/reg_to_wr_WB_reg[2]  ( .ip(n10068), .ck(clk), .q(
        \pipeline/reg_to_wr_WB [2]) );
  dp_1 \pipeline/ctrl/reg_to_wr_WB_reg[3]  ( .ip(n10067), .ck(clk), .q(
        \pipeline/reg_to_wr_WB [3]) );
  dp_1 \pipeline/dmem_type_WB_reg[0]  ( .ip(n8775), .ck(clk), .q(
        \pipeline/dmem_type_WB [0]) );
  dp_1 \pipeline/dmem_type_WB_reg[1]  ( .ip(n8774), .ck(clk), .q(
        \pipeline/dmem_type_WB [1]) );
  dp_1 \pipeline/dmem_type_WB_reg[2]  ( .ip(n8773), .ck(clk), .q(
        \pipeline/dmem_type_WB [2]) );
  dp_1 \pipeline/regfile/data_reg[1][0]  ( .ip(n9896), .ck(clk), .q(
        \pipeline/regfile/data[1][0] ) );
  dp_1 \pipeline/regfile/data_reg[1][1]  ( .ip(n9895), .ck(clk), .q(
        \pipeline/regfile/data[1][1] ) );
  dp_1 \pipeline/regfile/data_reg[1][2]  ( .ip(n9894), .ck(clk), .q(
        \pipeline/regfile/data[1][2] ) );
  dp_1 \pipeline/regfile/data_reg[1][3]  ( .ip(n9893), .ck(clk), .q(
        \pipeline/regfile/data[1][3] ) );
  dp_1 \pipeline/regfile/data_reg[1][4]  ( .ip(n9892), .ck(clk), .q(
        \pipeline/regfile/data[1][4] ) );
  dp_1 \pipeline/regfile/data_reg[1][5]  ( .ip(n9891), .ck(clk), .q(
        \pipeline/regfile/data[1][5] ) );
  dp_1 \pipeline/regfile/data_reg[1][6]  ( .ip(n9890), .ck(clk), .q(
        \pipeline/regfile/data[1][6] ) );
  dp_1 \pipeline/regfile/data_reg[1][7]  ( .ip(n9889), .ck(clk), .q(
        \pipeline/regfile/data[1][7] ) );
  dp_1 \pipeline/regfile/data_reg[1][8]  ( .ip(n9888), .ck(clk), .q(
        \pipeline/regfile/data[1][8] ) );
  dp_1 \pipeline/regfile/data_reg[1][9]  ( .ip(n9887), .ck(clk), .q(
        \pipeline/regfile/data[1][9] ) );
  dp_1 \pipeline/regfile/data_reg[1][10]  ( .ip(n9886), .ck(clk), .q(
        \pipeline/regfile/data[1][10] ) );
  dp_1 \pipeline/regfile/data_reg[1][11]  ( .ip(n9885), .ck(clk), .q(
        \pipeline/regfile/data[1][11] ) );
  dp_1 \pipeline/regfile/data_reg[1][12]  ( .ip(n9884), .ck(clk), .q(
        \pipeline/regfile/data[1][12] ) );
  dp_1 \pipeline/regfile/data_reg[1][13]  ( .ip(n9883), .ck(clk), .q(
        \pipeline/regfile/data[1][13] ) );
  dp_1 \pipeline/regfile/data_reg[1][14]  ( .ip(n9882), .ck(clk), .q(
        \pipeline/regfile/data[1][14] ) );
  dp_1 \pipeline/regfile/data_reg[1][15]  ( .ip(n9881), .ck(clk), .q(
        \pipeline/regfile/data[1][15] ) );
  dp_1 \pipeline/regfile/data_reg[1][16]  ( .ip(n9880), .ck(clk), .q(
        \pipeline/regfile/data[1][16] ) );
  dp_1 \pipeline/regfile/data_reg[1][17]  ( .ip(n9879), .ck(clk), .q(
        \pipeline/regfile/data[1][17] ) );
  dp_1 \pipeline/regfile/data_reg[1][18]  ( .ip(n9878), .ck(clk), .q(
        \pipeline/regfile/data[1][18] ) );
  dp_1 \pipeline/regfile/data_reg[1][19]  ( .ip(n9877), .ck(clk), .q(
        \pipeline/regfile/data[1][19] ) );
  dp_1 \pipeline/regfile/data_reg[1][20]  ( .ip(n9876), .ck(clk), .q(
        \pipeline/regfile/data[1][20] ) );
  dp_1 \pipeline/regfile/data_reg[1][21]  ( .ip(n9875), .ck(clk), .q(
        \pipeline/regfile/data[1][21] ) );
  dp_1 \pipeline/regfile/data_reg[1][22]  ( .ip(n9874), .ck(clk), .q(
        \pipeline/regfile/data[1][22] ) );
  dp_1 \pipeline/regfile/data_reg[1][23]  ( .ip(n9873), .ck(clk), .q(
        \pipeline/regfile/data[1][23] ) );
  dp_1 \pipeline/regfile/data_reg[1][24]  ( .ip(n9872), .ck(clk), .q(
        \pipeline/regfile/data[1][24] ) );
  dp_1 \pipeline/regfile/data_reg[1][25]  ( .ip(n9871), .ck(clk), .q(
        \pipeline/regfile/data[1][25] ) );
  dp_1 \pipeline/regfile/data_reg[1][26]  ( .ip(n9870), .ck(clk), .q(
        \pipeline/regfile/data[1][26] ) );
  dp_1 \pipeline/regfile/data_reg[1][27]  ( .ip(n9869), .ck(clk), .q(
        \pipeline/regfile/data[1][27] ) );
  dp_1 \pipeline/regfile/data_reg[1][28]  ( .ip(n9868), .ck(clk), .q(
        \pipeline/regfile/data[1][28] ) );
  dp_1 \pipeline/regfile/data_reg[1][29]  ( .ip(n9867), .ck(clk), .q(
        \pipeline/regfile/data[1][29] ) );
  dp_1 \pipeline/regfile/data_reg[1][30]  ( .ip(n9866), .ck(clk), .q(
        \pipeline/regfile/data[1][30] ) );
  dp_1 \pipeline/regfile/data_reg[1][31]  ( .ip(n9865), .ck(clk), .q(
        \pipeline/regfile/data[1][31] ) );
  dp_1 \pipeline/regfile/data_reg[2][0]  ( .ip(n9864), .ck(clk), .q(
        \pipeline/regfile/data[2][0] ) );
  dp_1 \pipeline/regfile/data_reg[2][1]  ( .ip(n9863), .ck(clk), .q(
        \pipeline/regfile/data[2][1] ) );
  dp_1 \pipeline/regfile/data_reg[2][2]  ( .ip(n9862), .ck(clk), .q(
        \pipeline/regfile/data[2][2] ) );
  dp_1 \pipeline/regfile/data_reg[2][3]  ( .ip(n9861), .ck(clk), .q(
        \pipeline/regfile/data[2][3] ) );
  dp_1 \pipeline/regfile/data_reg[2][4]  ( .ip(n9860), .ck(clk), .q(
        \pipeline/regfile/data[2][4] ) );
  dp_1 \pipeline/regfile/data_reg[2][5]  ( .ip(n9859), .ck(clk), .q(
        \pipeline/regfile/data[2][5] ) );
  dp_1 \pipeline/regfile/data_reg[2][6]  ( .ip(n9858), .ck(clk), .q(
        \pipeline/regfile/data[2][6] ) );
  dp_1 \pipeline/regfile/data_reg[2][7]  ( .ip(n9857), .ck(clk), .q(
        \pipeline/regfile/data[2][7] ) );
  dp_1 \pipeline/regfile/data_reg[2][8]  ( .ip(n9856), .ck(clk), .q(
        \pipeline/regfile/data[2][8] ) );
  dp_1 \pipeline/regfile/data_reg[2][9]  ( .ip(n9855), .ck(clk), .q(
        \pipeline/regfile/data[2][9] ) );
  dp_1 \pipeline/regfile/data_reg[2][10]  ( .ip(n9854), .ck(clk), .q(
        \pipeline/regfile/data[2][10] ) );
  dp_1 \pipeline/regfile/data_reg[2][11]  ( .ip(n9853), .ck(clk), .q(
        \pipeline/regfile/data[2][11] ) );
  dp_1 \pipeline/regfile/data_reg[2][12]  ( .ip(n9852), .ck(clk), .q(
        \pipeline/regfile/data[2][12] ) );
  dp_1 \pipeline/regfile/data_reg[2][13]  ( .ip(n9851), .ck(clk), .q(
        \pipeline/regfile/data[2][13] ) );
  dp_1 \pipeline/regfile/data_reg[2][14]  ( .ip(n9850), .ck(clk), .q(
        \pipeline/regfile/data[2][14] ) );
  dp_1 \pipeline/regfile/data_reg[2][15]  ( .ip(n9849), .ck(clk), .q(
        \pipeline/regfile/data[2][15] ) );
  dp_1 \pipeline/regfile/data_reg[2][16]  ( .ip(n9848), .ck(clk), .q(
        \pipeline/regfile/data[2][16] ) );
  dp_1 \pipeline/regfile/data_reg[2][17]  ( .ip(n9847), .ck(clk), .q(
        \pipeline/regfile/data[2][17] ) );
  dp_1 \pipeline/regfile/data_reg[2][18]  ( .ip(n9846), .ck(clk), .q(
        \pipeline/regfile/data[2][18] ) );
  dp_1 \pipeline/regfile/data_reg[2][19]  ( .ip(n9845), .ck(clk), .q(
        \pipeline/regfile/data[2][19] ) );
  dp_1 \pipeline/regfile/data_reg[2][20]  ( .ip(n9844), .ck(clk), .q(
        \pipeline/regfile/data[2][20] ) );
  dp_1 \pipeline/regfile/data_reg[2][21]  ( .ip(n9843), .ck(clk), .q(
        \pipeline/regfile/data[2][21] ) );
  dp_1 \pipeline/regfile/data_reg[2][22]  ( .ip(n9842), .ck(clk), .q(
        \pipeline/regfile/data[2][22] ) );
  dp_1 \pipeline/regfile/data_reg[2][23]  ( .ip(n9841), .ck(clk), .q(
        \pipeline/regfile/data[2][23] ) );
  dp_1 \pipeline/regfile/data_reg[2][24]  ( .ip(n9840), .ck(clk), .q(
        \pipeline/regfile/data[2][24] ) );
  dp_1 \pipeline/regfile/data_reg[2][25]  ( .ip(n9839), .ck(clk), .q(
        \pipeline/regfile/data[2][25] ) );
  dp_1 \pipeline/regfile/data_reg[2][26]  ( .ip(n9838), .ck(clk), .q(
        \pipeline/regfile/data[2][26] ) );
  dp_1 \pipeline/regfile/data_reg[2][27]  ( .ip(n9837), .ck(clk), .q(
        \pipeline/regfile/data[2][27] ) );
  dp_1 \pipeline/regfile/data_reg[2][28]  ( .ip(n9836), .ck(clk), .q(
        \pipeline/regfile/data[2][28] ) );
  dp_1 \pipeline/regfile/data_reg[2][29]  ( .ip(n9835), .ck(clk), .q(
        \pipeline/regfile/data[2][29] ) );
  dp_1 \pipeline/regfile/data_reg[2][30]  ( .ip(n9834), .ck(clk), .q(
        \pipeline/regfile/data[2][30] ) );
  dp_1 \pipeline/regfile/data_reg[2][31]  ( .ip(n9833), .ck(clk), .q(
        \pipeline/regfile/data[2][31] ) );
  dp_1 \pipeline/regfile/data_reg[3][0]  ( .ip(n9832), .ck(clk), .q(
        \pipeline/regfile/data[3][0] ) );
  dp_1 \pipeline/regfile/data_reg[3][1]  ( .ip(n9831), .ck(clk), .q(
        \pipeline/regfile/data[3][1] ) );
  dp_1 \pipeline/regfile/data_reg[3][2]  ( .ip(n9830), .ck(clk), .q(
        \pipeline/regfile/data[3][2] ) );
  dp_1 \pipeline/regfile/data_reg[3][3]  ( .ip(n9829), .ck(clk), .q(
        \pipeline/regfile/data[3][3] ) );
  dp_1 \pipeline/regfile/data_reg[3][4]  ( .ip(n9828), .ck(clk), .q(
        \pipeline/regfile/data[3][4] ) );
  dp_1 \pipeline/regfile/data_reg[3][5]  ( .ip(n9827), .ck(clk), .q(
        \pipeline/regfile/data[3][5] ) );
  dp_1 \pipeline/regfile/data_reg[3][6]  ( .ip(n9826), .ck(clk), .q(
        \pipeline/regfile/data[3][6] ) );
  dp_1 \pipeline/regfile/data_reg[3][7]  ( .ip(n9825), .ck(clk), .q(
        \pipeline/regfile/data[3][7] ) );
  dp_1 \pipeline/regfile/data_reg[3][8]  ( .ip(n9824), .ck(clk), .q(
        \pipeline/regfile/data[3][8] ) );
  dp_1 \pipeline/regfile/data_reg[3][9]  ( .ip(n9823), .ck(clk), .q(
        \pipeline/regfile/data[3][9] ) );
  dp_1 \pipeline/regfile/data_reg[3][10]  ( .ip(n9822), .ck(clk), .q(
        \pipeline/regfile/data[3][10] ) );
  dp_1 \pipeline/regfile/data_reg[3][11]  ( .ip(n9821), .ck(clk), .q(
        \pipeline/regfile/data[3][11] ) );
  dp_1 \pipeline/regfile/data_reg[3][12]  ( .ip(n9820), .ck(clk), .q(
        \pipeline/regfile/data[3][12] ) );
  dp_1 \pipeline/regfile/data_reg[3][13]  ( .ip(n9819), .ck(clk), .q(
        \pipeline/regfile/data[3][13] ) );
  dp_1 \pipeline/regfile/data_reg[3][14]  ( .ip(n9818), .ck(clk), .q(
        \pipeline/regfile/data[3][14] ) );
  dp_1 \pipeline/regfile/data_reg[3][15]  ( .ip(n9817), .ck(clk), .q(
        \pipeline/regfile/data[3][15] ) );
  dp_1 \pipeline/regfile/data_reg[3][16]  ( .ip(n9816), .ck(clk), .q(
        \pipeline/regfile/data[3][16] ) );
  dp_1 \pipeline/regfile/data_reg[3][17]  ( .ip(n9815), .ck(clk), .q(
        \pipeline/regfile/data[3][17] ) );
  dp_1 \pipeline/regfile/data_reg[3][18]  ( .ip(n9814), .ck(clk), .q(
        \pipeline/regfile/data[3][18] ) );
  dp_1 \pipeline/regfile/data_reg[3][19]  ( .ip(n9813), .ck(clk), .q(
        \pipeline/regfile/data[3][19] ) );
  dp_1 \pipeline/regfile/data_reg[3][20]  ( .ip(n9812), .ck(clk), .q(
        \pipeline/regfile/data[3][20] ) );
  dp_1 \pipeline/regfile/data_reg[3][21]  ( .ip(n9811), .ck(clk), .q(
        \pipeline/regfile/data[3][21] ) );
  dp_1 \pipeline/regfile/data_reg[3][22]  ( .ip(n9810), .ck(clk), .q(
        \pipeline/regfile/data[3][22] ) );
  dp_1 \pipeline/regfile/data_reg[3][23]  ( .ip(n9809), .ck(clk), .q(
        \pipeline/regfile/data[3][23] ) );
  dp_1 \pipeline/regfile/data_reg[3][24]  ( .ip(n9808), .ck(clk), .q(
        \pipeline/regfile/data[3][24] ) );
  dp_1 \pipeline/regfile/data_reg[3][25]  ( .ip(n9807), .ck(clk), .q(
        \pipeline/regfile/data[3][25] ) );
  dp_1 \pipeline/regfile/data_reg[3][26]  ( .ip(n9806), .ck(clk), .q(
        \pipeline/regfile/data[3][26] ) );
  dp_1 \pipeline/regfile/data_reg[3][27]  ( .ip(n9805), .ck(clk), .q(
        \pipeline/regfile/data[3][27] ) );
  dp_1 \pipeline/regfile/data_reg[3][28]  ( .ip(n9804), .ck(clk), .q(
        \pipeline/regfile/data[3][28] ) );
  dp_1 \pipeline/regfile/data_reg[3][29]  ( .ip(n9803), .ck(clk), .q(
        \pipeline/regfile/data[3][29] ) );
  dp_1 \pipeline/regfile/data_reg[3][30]  ( .ip(n9802), .ck(clk), .q(
        \pipeline/regfile/data[3][30] ) );
  dp_1 \pipeline/regfile/data_reg[3][31]  ( .ip(n9801), .ck(clk), .q(
        \pipeline/regfile/data[3][31] ) );
  dp_1 \pipeline/regfile/data_reg[4][0]  ( .ip(n9800), .ck(clk), .q(
        \pipeline/regfile/data[4][0] ) );
  dp_1 \pipeline/regfile/data_reg[4][1]  ( .ip(n9799), .ck(clk), .q(
        \pipeline/regfile/data[4][1] ) );
  dp_1 \pipeline/regfile/data_reg[4][2]  ( .ip(n9798), .ck(clk), .q(
        \pipeline/regfile/data[4][2] ) );
  dp_1 \pipeline/regfile/data_reg[4][3]  ( .ip(n9797), .ck(clk), .q(
        \pipeline/regfile/data[4][3] ) );
  dp_1 \pipeline/regfile/data_reg[4][4]  ( .ip(n9796), .ck(clk), .q(
        \pipeline/regfile/data[4][4] ) );
  dp_1 \pipeline/regfile/data_reg[4][5]  ( .ip(n9795), .ck(clk), .q(
        \pipeline/regfile/data[4][5] ) );
  dp_1 \pipeline/regfile/data_reg[4][6]  ( .ip(n9794), .ck(clk), .q(
        \pipeline/regfile/data[4][6] ) );
  dp_1 \pipeline/regfile/data_reg[4][7]  ( .ip(n9793), .ck(clk), .q(
        \pipeline/regfile/data[4][7] ) );
  dp_1 \pipeline/regfile/data_reg[4][8]  ( .ip(n9792), .ck(clk), .q(
        \pipeline/regfile/data[4][8] ) );
  dp_1 \pipeline/regfile/data_reg[4][9]  ( .ip(n9791), .ck(clk), .q(
        \pipeline/regfile/data[4][9] ) );
  dp_1 \pipeline/regfile/data_reg[4][10]  ( .ip(n9790), .ck(clk), .q(
        \pipeline/regfile/data[4][10] ) );
  dp_1 \pipeline/regfile/data_reg[4][11]  ( .ip(n9789), .ck(clk), .q(
        \pipeline/regfile/data[4][11] ) );
  dp_1 \pipeline/regfile/data_reg[4][12]  ( .ip(n9788), .ck(clk), .q(
        \pipeline/regfile/data[4][12] ) );
  dp_1 \pipeline/regfile/data_reg[4][13]  ( .ip(n9787), .ck(clk), .q(
        \pipeline/regfile/data[4][13] ) );
  dp_1 \pipeline/regfile/data_reg[4][14]  ( .ip(n9786), .ck(clk), .q(
        \pipeline/regfile/data[4][14] ) );
  dp_1 \pipeline/regfile/data_reg[4][15]  ( .ip(n9785), .ck(clk), .q(
        \pipeline/regfile/data[4][15] ) );
  dp_1 \pipeline/regfile/data_reg[4][16]  ( .ip(n9784), .ck(clk), .q(
        \pipeline/regfile/data[4][16] ) );
  dp_1 \pipeline/regfile/data_reg[4][17]  ( .ip(n9783), .ck(clk), .q(
        \pipeline/regfile/data[4][17] ) );
  dp_1 \pipeline/regfile/data_reg[4][18]  ( .ip(n9782), .ck(clk), .q(
        \pipeline/regfile/data[4][18] ) );
  dp_1 \pipeline/regfile/data_reg[4][19]  ( .ip(n9781), .ck(clk), .q(
        \pipeline/regfile/data[4][19] ) );
  dp_1 \pipeline/regfile/data_reg[4][20]  ( .ip(n9780), .ck(clk), .q(
        \pipeline/regfile/data[4][20] ) );
  dp_1 \pipeline/regfile/data_reg[4][21]  ( .ip(n9779), .ck(clk), .q(
        \pipeline/regfile/data[4][21] ) );
  dp_1 \pipeline/regfile/data_reg[4][22]  ( .ip(n9778), .ck(clk), .q(
        \pipeline/regfile/data[4][22] ) );
  dp_1 \pipeline/regfile/data_reg[4][23]  ( .ip(n9777), .ck(clk), .q(
        \pipeline/regfile/data[4][23] ) );
  dp_1 \pipeline/regfile/data_reg[4][24]  ( .ip(n9776), .ck(clk), .q(
        \pipeline/regfile/data[4][24] ) );
  dp_1 \pipeline/regfile/data_reg[4][25]  ( .ip(n9775), .ck(clk), .q(
        \pipeline/regfile/data[4][25] ) );
  dp_1 \pipeline/regfile/data_reg[4][26]  ( .ip(n9774), .ck(clk), .q(
        \pipeline/regfile/data[4][26] ) );
  dp_1 \pipeline/regfile/data_reg[4][27]  ( .ip(n9773), .ck(clk), .q(
        \pipeline/regfile/data[4][27] ) );
  dp_1 \pipeline/regfile/data_reg[4][28]  ( .ip(n9772), .ck(clk), .q(
        \pipeline/regfile/data[4][28] ) );
  dp_1 \pipeline/regfile/data_reg[4][29]  ( .ip(n9771), .ck(clk), .q(
        \pipeline/regfile/data[4][29] ) );
  dp_1 \pipeline/regfile/data_reg[4][30]  ( .ip(n9770), .ck(clk), .q(
        \pipeline/regfile/data[4][30] ) );
  dp_1 \pipeline/regfile/data_reg[4][31]  ( .ip(n9769), .ck(clk), .q(
        \pipeline/regfile/data[4][31] ) );
  dp_1 \pipeline/regfile/data_reg[5][0]  ( .ip(n9768), .ck(clk), .q(
        \pipeline/regfile/data[5][0] ) );
  dp_1 \pipeline/regfile/data_reg[5][1]  ( .ip(n9767), .ck(clk), .q(
        \pipeline/regfile/data[5][1] ) );
  dp_1 \pipeline/regfile/data_reg[5][2]  ( .ip(n9766), .ck(clk), .q(
        \pipeline/regfile/data[5][2] ) );
  dp_1 \pipeline/regfile/data_reg[5][3]  ( .ip(n9765), .ck(clk), .q(
        \pipeline/regfile/data[5][3] ) );
  dp_1 \pipeline/regfile/data_reg[5][4]  ( .ip(n9764), .ck(clk), .q(
        \pipeline/regfile/data[5][4] ) );
  dp_1 \pipeline/regfile/data_reg[5][5]  ( .ip(n9763), .ck(clk), .q(
        \pipeline/regfile/data[5][5] ) );
  dp_1 \pipeline/regfile/data_reg[5][6]  ( .ip(n9762), .ck(clk), .q(
        \pipeline/regfile/data[5][6] ) );
  dp_1 \pipeline/regfile/data_reg[5][7]  ( .ip(n9761), .ck(clk), .q(
        \pipeline/regfile/data[5][7] ) );
  dp_1 \pipeline/regfile/data_reg[5][8]  ( .ip(n9760), .ck(clk), .q(
        \pipeline/regfile/data[5][8] ) );
  dp_1 \pipeline/regfile/data_reg[5][9]  ( .ip(n9759), .ck(clk), .q(
        \pipeline/regfile/data[5][9] ) );
  dp_1 \pipeline/regfile/data_reg[5][10]  ( .ip(n9758), .ck(clk), .q(
        \pipeline/regfile/data[5][10] ) );
  dp_1 \pipeline/regfile/data_reg[5][11]  ( .ip(n9757), .ck(clk), .q(
        \pipeline/regfile/data[5][11] ) );
  dp_1 \pipeline/regfile/data_reg[5][12]  ( .ip(n9756), .ck(clk), .q(
        \pipeline/regfile/data[5][12] ) );
  dp_1 \pipeline/regfile/data_reg[5][13]  ( .ip(n9755), .ck(clk), .q(
        \pipeline/regfile/data[5][13] ) );
  dp_1 \pipeline/regfile/data_reg[5][14]  ( .ip(n9754), .ck(clk), .q(
        \pipeline/regfile/data[5][14] ) );
  dp_1 \pipeline/regfile/data_reg[5][15]  ( .ip(n9753), .ck(clk), .q(
        \pipeline/regfile/data[5][15] ) );
  dp_1 \pipeline/regfile/data_reg[5][16]  ( .ip(n9752), .ck(clk), .q(
        \pipeline/regfile/data[5][16] ) );
  dp_1 \pipeline/regfile/data_reg[5][17]  ( .ip(n9751), .ck(clk), .q(
        \pipeline/regfile/data[5][17] ) );
  dp_1 \pipeline/regfile/data_reg[5][18]  ( .ip(n9750), .ck(clk), .q(
        \pipeline/regfile/data[5][18] ) );
  dp_1 \pipeline/regfile/data_reg[5][19]  ( .ip(n9749), .ck(clk), .q(
        \pipeline/regfile/data[5][19] ) );
  dp_1 \pipeline/regfile/data_reg[5][20]  ( .ip(n9748), .ck(clk), .q(
        \pipeline/regfile/data[5][20] ) );
  dp_1 \pipeline/regfile/data_reg[5][21]  ( .ip(n9747), .ck(clk), .q(
        \pipeline/regfile/data[5][21] ) );
  dp_1 \pipeline/regfile/data_reg[5][22]  ( .ip(n9746), .ck(clk), .q(
        \pipeline/regfile/data[5][22] ) );
  dp_1 \pipeline/regfile/data_reg[5][23]  ( .ip(n9745), .ck(clk), .q(
        \pipeline/regfile/data[5][23] ) );
  dp_1 \pipeline/regfile/data_reg[5][24]  ( .ip(n9744), .ck(clk), .q(
        \pipeline/regfile/data[5][24] ) );
  dp_1 \pipeline/regfile/data_reg[5][25]  ( .ip(n9743), .ck(clk), .q(
        \pipeline/regfile/data[5][25] ) );
  dp_1 \pipeline/regfile/data_reg[5][26]  ( .ip(n9742), .ck(clk), .q(
        \pipeline/regfile/data[5][26] ) );
  dp_1 \pipeline/regfile/data_reg[5][27]  ( .ip(n9741), .ck(clk), .q(
        \pipeline/regfile/data[5][27] ) );
  dp_1 \pipeline/regfile/data_reg[5][28]  ( .ip(n9740), .ck(clk), .q(
        \pipeline/regfile/data[5][28] ) );
  dp_1 \pipeline/regfile/data_reg[5][29]  ( .ip(n9739), .ck(clk), .q(
        \pipeline/regfile/data[5][29] ) );
  dp_1 \pipeline/regfile/data_reg[5][30]  ( .ip(n9738), .ck(clk), .q(
        \pipeline/regfile/data[5][30] ) );
  dp_1 \pipeline/regfile/data_reg[5][31]  ( .ip(n9737), .ck(clk), .q(
        \pipeline/regfile/data[5][31] ) );
  dp_1 \pipeline/regfile/data_reg[6][0]  ( .ip(n9736), .ck(clk), .q(
        \pipeline/regfile/data[6][0] ) );
  dp_1 \pipeline/regfile/data_reg[6][1]  ( .ip(n9735), .ck(clk), .q(
        \pipeline/regfile/data[6][1] ) );
  dp_1 \pipeline/regfile/data_reg[6][2]  ( .ip(n9734), .ck(clk), .q(
        \pipeline/regfile/data[6][2] ) );
  dp_1 \pipeline/regfile/data_reg[6][3]  ( .ip(n9733), .ck(clk), .q(
        \pipeline/regfile/data[6][3] ) );
  dp_1 \pipeline/regfile/data_reg[6][4]  ( .ip(n9732), .ck(clk), .q(
        \pipeline/regfile/data[6][4] ) );
  dp_1 \pipeline/regfile/data_reg[6][5]  ( .ip(n9731), .ck(clk), .q(
        \pipeline/regfile/data[6][5] ) );
  dp_1 \pipeline/regfile/data_reg[6][6]  ( .ip(n9730), .ck(clk), .q(
        \pipeline/regfile/data[6][6] ) );
  dp_1 \pipeline/regfile/data_reg[6][7]  ( .ip(n9729), .ck(clk), .q(
        \pipeline/regfile/data[6][7] ) );
  dp_1 \pipeline/regfile/data_reg[6][8]  ( .ip(n9728), .ck(clk), .q(
        \pipeline/regfile/data[6][8] ) );
  dp_1 \pipeline/regfile/data_reg[6][9]  ( .ip(n9727), .ck(clk), .q(
        \pipeline/regfile/data[6][9] ) );
  dp_1 \pipeline/regfile/data_reg[6][10]  ( .ip(n9726), .ck(clk), .q(
        \pipeline/regfile/data[6][10] ) );
  dp_1 \pipeline/regfile/data_reg[6][11]  ( .ip(n9725), .ck(clk), .q(
        \pipeline/regfile/data[6][11] ) );
  dp_1 \pipeline/regfile/data_reg[6][12]  ( .ip(n9724), .ck(clk), .q(
        \pipeline/regfile/data[6][12] ) );
  dp_1 \pipeline/regfile/data_reg[6][13]  ( .ip(n9723), .ck(clk), .q(
        \pipeline/regfile/data[6][13] ) );
  dp_1 \pipeline/regfile/data_reg[6][14]  ( .ip(n9722), .ck(clk), .q(
        \pipeline/regfile/data[6][14] ) );
  dp_1 \pipeline/regfile/data_reg[6][15]  ( .ip(n9721), .ck(clk), .q(
        \pipeline/regfile/data[6][15] ) );
  dp_1 \pipeline/regfile/data_reg[6][16]  ( .ip(n9720), .ck(clk), .q(
        \pipeline/regfile/data[6][16] ) );
  dp_1 \pipeline/regfile/data_reg[6][17]  ( .ip(n9719), .ck(clk), .q(
        \pipeline/regfile/data[6][17] ) );
  dp_1 \pipeline/regfile/data_reg[6][18]  ( .ip(n9718), .ck(clk), .q(
        \pipeline/regfile/data[6][18] ) );
  dp_1 \pipeline/regfile/data_reg[6][19]  ( .ip(n9717), .ck(clk), .q(
        \pipeline/regfile/data[6][19] ) );
  dp_1 \pipeline/regfile/data_reg[6][20]  ( .ip(n9716), .ck(clk), .q(
        \pipeline/regfile/data[6][20] ) );
  dp_1 \pipeline/regfile/data_reg[6][21]  ( .ip(n9715), .ck(clk), .q(
        \pipeline/regfile/data[6][21] ) );
  dp_1 \pipeline/regfile/data_reg[6][22]  ( .ip(n9714), .ck(clk), .q(
        \pipeline/regfile/data[6][22] ) );
  dp_1 \pipeline/regfile/data_reg[6][23]  ( .ip(n9713), .ck(clk), .q(
        \pipeline/regfile/data[6][23] ) );
  dp_1 \pipeline/regfile/data_reg[6][24]  ( .ip(n9712), .ck(clk), .q(
        \pipeline/regfile/data[6][24] ) );
  dp_1 \pipeline/regfile/data_reg[6][25]  ( .ip(n9711), .ck(clk), .q(
        \pipeline/regfile/data[6][25] ) );
  dp_1 \pipeline/regfile/data_reg[6][26]  ( .ip(n9710), .ck(clk), .q(
        \pipeline/regfile/data[6][26] ) );
  dp_1 \pipeline/regfile/data_reg[6][27]  ( .ip(n9709), .ck(clk), .q(
        \pipeline/regfile/data[6][27] ) );
  dp_1 \pipeline/regfile/data_reg[6][28]  ( .ip(n9708), .ck(clk), .q(
        \pipeline/regfile/data[6][28] ) );
  dp_1 \pipeline/regfile/data_reg[6][29]  ( .ip(n9707), .ck(clk), .q(
        \pipeline/regfile/data[6][29] ) );
  dp_1 \pipeline/regfile/data_reg[6][30]  ( .ip(n9706), .ck(clk), .q(
        \pipeline/regfile/data[6][30] ) );
  dp_1 \pipeline/regfile/data_reg[6][31]  ( .ip(n9705), .ck(clk), .q(
        \pipeline/regfile/data[6][31] ) );
  dp_1 \pipeline/regfile/data_reg[7][0]  ( .ip(n9704), .ck(clk), .q(
        \pipeline/regfile/data[7][0] ) );
  dp_1 \pipeline/regfile/data_reg[7][1]  ( .ip(n9703), .ck(clk), .q(
        \pipeline/regfile/data[7][1] ) );
  dp_1 \pipeline/regfile/data_reg[7][2]  ( .ip(n9702), .ck(clk), .q(
        \pipeline/regfile/data[7][2] ) );
  dp_1 \pipeline/regfile/data_reg[7][3]  ( .ip(n9701), .ck(clk), .q(
        \pipeline/regfile/data[7][3] ) );
  dp_1 \pipeline/regfile/data_reg[7][4]  ( .ip(n9700), .ck(clk), .q(
        \pipeline/regfile/data[7][4] ) );
  dp_1 \pipeline/regfile/data_reg[7][5]  ( .ip(n9699), .ck(clk), .q(
        \pipeline/regfile/data[7][5] ) );
  dp_1 \pipeline/regfile/data_reg[7][6]  ( .ip(n9698), .ck(clk), .q(
        \pipeline/regfile/data[7][6] ) );
  dp_1 \pipeline/regfile/data_reg[7][7]  ( .ip(n9697), .ck(clk), .q(
        \pipeline/regfile/data[7][7] ) );
  dp_1 \pipeline/regfile/data_reg[7][8]  ( .ip(n9696), .ck(clk), .q(
        \pipeline/regfile/data[7][8] ) );
  dp_1 \pipeline/regfile/data_reg[7][9]  ( .ip(n9695), .ck(clk), .q(
        \pipeline/regfile/data[7][9] ) );
  dp_1 \pipeline/regfile/data_reg[7][10]  ( .ip(n9694), .ck(clk), .q(
        \pipeline/regfile/data[7][10] ) );
  dp_1 \pipeline/regfile/data_reg[7][11]  ( .ip(n9693), .ck(clk), .q(
        \pipeline/regfile/data[7][11] ) );
  dp_1 \pipeline/regfile/data_reg[7][12]  ( .ip(n9692), .ck(clk), .q(
        \pipeline/regfile/data[7][12] ) );
  dp_1 \pipeline/regfile/data_reg[7][13]  ( .ip(n9691), .ck(clk), .q(
        \pipeline/regfile/data[7][13] ) );
  dp_1 \pipeline/regfile/data_reg[7][14]  ( .ip(n9690), .ck(clk), .q(
        \pipeline/regfile/data[7][14] ) );
  dp_1 \pipeline/regfile/data_reg[7][15]  ( .ip(n9689), .ck(clk), .q(
        \pipeline/regfile/data[7][15] ) );
  dp_1 \pipeline/regfile/data_reg[7][16]  ( .ip(n9688), .ck(clk), .q(
        \pipeline/regfile/data[7][16] ) );
  dp_1 \pipeline/regfile/data_reg[7][17]  ( .ip(n9687), .ck(clk), .q(
        \pipeline/regfile/data[7][17] ) );
  dp_1 \pipeline/regfile/data_reg[7][18]  ( .ip(n9686), .ck(clk), .q(
        \pipeline/regfile/data[7][18] ) );
  dp_1 \pipeline/regfile/data_reg[7][19]  ( .ip(n9685), .ck(clk), .q(
        \pipeline/regfile/data[7][19] ) );
  dp_1 \pipeline/regfile/data_reg[7][20]  ( .ip(n9684), .ck(clk), .q(
        \pipeline/regfile/data[7][20] ) );
  dp_1 \pipeline/regfile/data_reg[7][21]  ( .ip(n9683), .ck(clk), .q(
        \pipeline/regfile/data[7][21] ) );
  dp_1 \pipeline/regfile/data_reg[7][22]  ( .ip(n9682), .ck(clk), .q(
        \pipeline/regfile/data[7][22] ) );
  dp_1 \pipeline/regfile/data_reg[7][23]  ( .ip(n9681), .ck(clk), .q(
        \pipeline/regfile/data[7][23] ) );
  dp_1 \pipeline/regfile/data_reg[7][24]  ( .ip(n9680), .ck(clk), .q(
        \pipeline/regfile/data[7][24] ) );
  dp_1 \pipeline/regfile/data_reg[7][25]  ( .ip(n9679), .ck(clk), .q(
        \pipeline/regfile/data[7][25] ) );
  dp_1 \pipeline/regfile/data_reg[7][26]  ( .ip(n9678), .ck(clk), .q(
        \pipeline/regfile/data[7][26] ) );
  dp_1 \pipeline/regfile/data_reg[7][27]  ( .ip(n9677), .ck(clk), .q(
        \pipeline/regfile/data[7][27] ) );
  dp_1 \pipeline/regfile/data_reg[7][28]  ( .ip(n9676), .ck(clk), .q(
        \pipeline/regfile/data[7][28] ) );
  dp_1 \pipeline/regfile/data_reg[7][29]  ( .ip(n9675), .ck(clk), .q(
        \pipeline/regfile/data[7][29] ) );
  dp_1 \pipeline/regfile/data_reg[7][30]  ( .ip(n9674), .ck(clk), .q(
        \pipeline/regfile/data[7][30] ) );
  dp_1 \pipeline/regfile/data_reg[7][31]  ( .ip(n9673), .ck(clk), .q(
        \pipeline/regfile/data[7][31] ) );
  dp_1 \pipeline/regfile/data_reg[8][0]  ( .ip(n9672), .ck(clk), .q(
        \pipeline/regfile/data[8][0] ) );
  dp_1 \pipeline/regfile/data_reg[8][1]  ( .ip(n9671), .ck(clk), .q(
        \pipeline/regfile/data[8][1] ) );
  dp_1 \pipeline/regfile/data_reg[8][2]  ( .ip(n9670), .ck(clk), .q(
        \pipeline/regfile/data[8][2] ) );
  dp_1 \pipeline/regfile/data_reg[8][3]  ( .ip(n9669), .ck(clk), .q(
        \pipeline/regfile/data[8][3] ) );
  dp_1 \pipeline/regfile/data_reg[8][4]  ( .ip(n9668), .ck(clk), .q(
        \pipeline/regfile/data[8][4] ) );
  dp_1 \pipeline/regfile/data_reg[8][5]  ( .ip(n9667), .ck(clk), .q(
        \pipeline/regfile/data[8][5] ) );
  dp_1 \pipeline/regfile/data_reg[8][6]  ( .ip(n9666), .ck(clk), .q(
        \pipeline/regfile/data[8][6] ) );
  dp_1 \pipeline/regfile/data_reg[8][7]  ( .ip(n9665), .ck(clk), .q(
        \pipeline/regfile/data[8][7] ) );
  dp_1 \pipeline/regfile/data_reg[8][8]  ( .ip(n9664), .ck(clk), .q(
        \pipeline/regfile/data[8][8] ) );
  dp_1 \pipeline/regfile/data_reg[8][9]  ( .ip(n9663), .ck(clk), .q(
        \pipeline/regfile/data[8][9] ) );
  dp_1 \pipeline/regfile/data_reg[8][10]  ( .ip(n9662), .ck(clk), .q(
        \pipeline/regfile/data[8][10] ) );
  dp_1 \pipeline/regfile/data_reg[8][11]  ( .ip(n9661), .ck(clk), .q(
        \pipeline/regfile/data[8][11] ) );
  dp_1 \pipeline/regfile/data_reg[8][12]  ( .ip(n9660), .ck(clk), .q(
        \pipeline/regfile/data[8][12] ) );
  dp_1 \pipeline/regfile/data_reg[8][13]  ( .ip(n9659), .ck(clk), .q(
        \pipeline/regfile/data[8][13] ) );
  dp_1 \pipeline/regfile/data_reg[8][14]  ( .ip(n9658), .ck(clk), .q(
        \pipeline/regfile/data[8][14] ) );
  dp_1 \pipeline/regfile/data_reg[8][15]  ( .ip(n9657), .ck(clk), .q(
        \pipeline/regfile/data[8][15] ) );
  dp_1 \pipeline/regfile/data_reg[8][16]  ( .ip(n9656), .ck(clk), .q(
        \pipeline/regfile/data[8][16] ) );
  dp_1 \pipeline/regfile/data_reg[8][17]  ( .ip(n9655), .ck(clk), .q(
        \pipeline/regfile/data[8][17] ) );
  dp_1 \pipeline/regfile/data_reg[8][18]  ( .ip(n9654), .ck(clk), .q(
        \pipeline/regfile/data[8][18] ) );
  dp_1 \pipeline/regfile/data_reg[8][19]  ( .ip(n9653), .ck(clk), .q(
        \pipeline/regfile/data[8][19] ) );
  dp_1 \pipeline/regfile/data_reg[8][20]  ( .ip(n9652), .ck(clk), .q(
        \pipeline/regfile/data[8][20] ) );
  dp_1 \pipeline/regfile/data_reg[8][21]  ( .ip(n9651), .ck(clk), .q(
        \pipeline/regfile/data[8][21] ) );
  dp_1 \pipeline/regfile/data_reg[8][22]  ( .ip(n9650), .ck(clk), .q(
        \pipeline/regfile/data[8][22] ) );
  dp_1 \pipeline/regfile/data_reg[8][23]  ( .ip(n9649), .ck(clk), .q(
        \pipeline/regfile/data[8][23] ) );
  dp_1 \pipeline/regfile/data_reg[8][24]  ( .ip(n9648), .ck(clk), .q(
        \pipeline/regfile/data[8][24] ) );
  dp_1 \pipeline/regfile/data_reg[8][25]  ( .ip(n9647), .ck(clk), .q(
        \pipeline/regfile/data[8][25] ) );
  dp_1 \pipeline/regfile/data_reg[8][26]  ( .ip(n9646), .ck(clk), .q(
        \pipeline/regfile/data[8][26] ) );
  dp_1 \pipeline/regfile/data_reg[8][27]  ( .ip(n9645), .ck(clk), .q(
        \pipeline/regfile/data[8][27] ) );
  dp_1 \pipeline/regfile/data_reg[8][28]  ( .ip(n9644), .ck(clk), .q(
        \pipeline/regfile/data[8][28] ) );
  dp_1 \pipeline/regfile/data_reg[8][29]  ( .ip(n9643), .ck(clk), .q(
        \pipeline/regfile/data[8][29] ) );
  dp_1 \pipeline/regfile/data_reg[8][30]  ( .ip(n9642), .ck(clk), .q(
        \pipeline/regfile/data[8][30] ) );
  dp_1 \pipeline/regfile/data_reg[8][31]  ( .ip(n9641), .ck(clk), .q(
        \pipeline/regfile/data[8][31] ) );
  dp_1 \pipeline/regfile/data_reg[9][0]  ( .ip(n9640), .ck(clk), .q(
        \pipeline/regfile/data[9][0] ) );
  dp_1 \pipeline/regfile/data_reg[9][1]  ( .ip(n9639), .ck(clk), .q(
        \pipeline/regfile/data[9][1] ) );
  dp_1 \pipeline/regfile/data_reg[9][2]  ( .ip(n9638), .ck(clk), .q(
        \pipeline/regfile/data[9][2] ) );
  dp_1 \pipeline/regfile/data_reg[9][3]  ( .ip(n9637), .ck(clk), .q(
        \pipeline/regfile/data[9][3] ) );
  dp_1 \pipeline/regfile/data_reg[9][4]  ( .ip(n9636), .ck(clk), .q(
        \pipeline/regfile/data[9][4] ) );
  dp_1 \pipeline/regfile/data_reg[9][5]  ( .ip(n9635), .ck(clk), .q(
        \pipeline/regfile/data[9][5] ) );
  dp_1 \pipeline/regfile/data_reg[9][6]  ( .ip(n9634), .ck(clk), .q(
        \pipeline/regfile/data[9][6] ) );
  dp_1 \pipeline/regfile/data_reg[9][7]  ( .ip(n9633), .ck(clk), .q(
        \pipeline/regfile/data[9][7] ) );
  dp_1 \pipeline/regfile/data_reg[9][8]  ( .ip(n9632), .ck(clk), .q(
        \pipeline/regfile/data[9][8] ) );
  dp_1 \pipeline/regfile/data_reg[9][9]  ( .ip(n9631), .ck(clk), .q(
        \pipeline/regfile/data[9][9] ) );
  dp_1 \pipeline/regfile/data_reg[9][10]  ( .ip(n9630), .ck(clk), .q(
        \pipeline/regfile/data[9][10] ) );
  dp_1 \pipeline/regfile/data_reg[9][11]  ( .ip(n9629), .ck(clk), .q(
        \pipeline/regfile/data[9][11] ) );
  dp_1 \pipeline/regfile/data_reg[9][12]  ( .ip(n9628), .ck(clk), .q(
        \pipeline/regfile/data[9][12] ) );
  dp_1 \pipeline/regfile/data_reg[9][13]  ( .ip(n9627), .ck(clk), .q(
        \pipeline/regfile/data[9][13] ) );
  dp_1 \pipeline/regfile/data_reg[9][14]  ( .ip(n9626), .ck(clk), .q(
        \pipeline/regfile/data[9][14] ) );
  dp_1 \pipeline/regfile/data_reg[9][15]  ( .ip(n9625), .ck(clk), .q(
        \pipeline/regfile/data[9][15] ) );
  dp_1 \pipeline/regfile/data_reg[9][16]  ( .ip(n9624), .ck(clk), .q(
        \pipeline/regfile/data[9][16] ) );
  dp_1 \pipeline/regfile/data_reg[9][17]  ( .ip(n9623), .ck(clk), .q(
        \pipeline/regfile/data[9][17] ) );
  dp_1 \pipeline/regfile/data_reg[9][18]  ( .ip(n9622), .ck(clk), .q(
        \pipeline/regfile/data[9][18] ) );
  dp_1 \pipeline/regfile/data_reg[9][19]  ( .ip(n9621), .ck(clk), .q(
        \pipeline/regfile/data[9][19] ) );
  dp_1 \pipeline/regfile/data_reg[9][20]  ( .ip(n9620), .ck(clk), .q(
        \pipeline/regfile/data[9][20] ) );
  dp_1 \pipeline/regfile/data_reg[9][21]  ( .ip(n9619), .ck(clk), .q(
        \pipeline/regfile/data[9][21] ) );
  dp_1 \pipeline/regfile/data_reg[9][22]  ( .ip(n9618), .ck(clk), .q(
        \pipeline/regfile/data[9][22] ) );
  dp_1 \pipeline/regfile/data_reg[9][23]  ( .ip(n9617), .ck(clk), .q(
        \pipeline/regfile/data[9][23] ) );
  dp_1 \pipeline/regfile/data_reg[9][24]  ( .ip(n9616), .ck(clk), .q(
        \pipeline/regfile/data[9][24] ) );
  dp_1 \pipeline/regfile/data_reg[9][25]  ( .ip(n9615), .ck(clk), .q(
        \pipeline/regfile/data[9][25] ) );
  dp_1 \pipeline/regfile/data_reg[9][26]  ( .ip(n9614), .ck(clk), .q(
        \pipeline/regfile/data[9][26] ) );
  dp_1 \pipeline/regfile/data_reg[9][27]  ( .ip(n9613), .ck(clk), .q(
        \pipeline/regfile/data[9][27] ) );
  dp_1 \pipeline/regfile/data_reg[9][28]  ( .ip(n9612), .ck(clk), .q(
        \pipeline/regfile/data[9][28] ) );
  dp_1 \pipeline/regfile/data_reg[9][29]  ( .ip(n9611), .ck(clk), .q(
        \pipeline/regfile/data[9][29] ) );
  dp_1 \pipeline/regfile/data_reg[9][30]  ( .ip(n9610), .ck(clk), .q(
        \pipeline/regfile/data[9][30] ) );
  dp_1 \pipeline/regfile/data_reg[9][31]  ( .ip(n9609), .ck(clk), .q(
        \pipeline/regfile/data[9][31] ) );
  dp_1 \pipeline/regfile/data_reg[10][0]  ( .ip(n9608), .ck(clk), .q(
        \pipeline/regfile/data[10][0] ) );
  dp_1 \pipeline/regfile/data_reg[10][1]  ( .ip(n9607), .ck(clk), .q(
        \pipeline/regfile/data[10][1] ) );
  dp_1 \pipeline/regfile/data_reg[10][2]  ( .ip(n9606), .ck(clk), .q(
        \pipeline/regfile/data[10][2] ) );
  dp_1 \pipeline/regfile/data_reg[10][3]  ( .ip(n9605), .ck(clk), .q(
        \pipeline/regfile/data[10][3] ) );
  dp_1 \pipeline/regfile/data_reg[10][4]  ( .ip(n9604), .ck(clk), .q(
        \pipeline/regfile/data[10][4] ) );
  dp_1 \pipeline/regfile/data_reg[10][5]  ( .ip(n9603), .ck(clk), .q(
        \pipeline/regfile/data[10][5] ) );
  dp_1 \pipeline/regfile/data_reg[10][6]  ( .ip(n9602), .ck(clk), .q(
        \pipeline/regfile/data[10][6] ) );
  dp_1 \pipeline/regfile/data_reg[10][7]  ( .ip(n9601), .ck(clk), .q(
        \pipeline/regfile/data[10][7] ) );
  dp_1 \pipeline/regfile/data_reg[10][8]  ( .ip(n9600), .ck(clk), .q(
        \pipeline/regfile/data[10][8] ) );
  dp_1 \pipeline/regfile/data_reg[10][9]  ( .ip(n9599), .ck(clk), .q(
        \pipeline/regfile/data[10][9] ) );
  dp_1 \pipeline/regfile/data_reg[10][10]  ( .ip(n9598), .ck(clk), .q(
        \pipeline/regfile/data[10][10] ) );
  dp_1 \pipeline/regfile/data_reg[10][11]  ( .ip(n9597), .ck(clk), .q(
        \pipeline/regfile/data[10][11] ) );
  dp_1 \pipeline/regfile/data_reg[10][12]  ( .ip(n9596), .ck(clk), .q(
        \pipeline/regfile/data[10][12] ) );
  dp_1 \pipeline/regfile/data_reg[10][13]  ( .ip(n9595), .ck(clk), .q(
        \pipeline/regfile/data[10][13] ) );
  dp_1 \pipeline/regfile/data_reg[10][14]  ( .ip(n9594), .ck(clk), .q(
        \pipeline/regfile/data[10][14] ) );
  dp_1 \pipeline/regfile/data_reg[10][15]  ( .ip(n9593), .ck(clk), .q(
        \pipeline/regfile/data[10][15] ) );
  dp_1 \pipeline/regfile/data_reg[10][16]  ( .ip(n9592), .ck(clk), .q(
        \pipeline/regfile/data[10][16] ) );
  dp_1 \pipeline/regfile/data_reg[10][17]  ( .ip(n9591), .ck(clk), .q(
        \pipeline/regfile/data[10][17] ) );
  dp_1 \pipeline/regfile/data_reg[10][18]  ( .ip(n9590), .ck(clk), .q(
        \pipeline/regfile/data[10][18] ) );
  dp_1 \pipeline/regfile/data_reg[10][19]  ( .ip(n9589), .ck(clk), .q(
        \pipeline/regfile/data[10][19] ) );
  dp_1 \pipeline/regfile/data_reg[10][20]  ( .ip(n9588), .ck(clk), .q(
        \pipeline/regfile/data[10][20] ) );
  dp_1 \pipeline/regfile/data_reg[10][21]  ( .ip(n9587), .ck(clk), .q(
        \pipeline/regfile/data[10][21] ) );
  dp_1 \pipeline/regfile/data_reg[10][22]  ( .ip(n9586), .ck(clk), .q(
        \pipeline/regfile/data[10][22] ) );
  dp_1 \pipeline/regfile/data_reg[10][23]  ( .ip(n9585), .ck(clk), .q(
        \pipeline/regfile/data[10][23] ) );
  dp_1 \pipeline/regfile/data_reg[10][24]  ( .ip(n9584), .ck(clk), .q(
        \pipeline/regfile/data[10][24] ) );
  dp_1 \pipeline/regfile/data_reg[10][25]  ( .ip(n9583), .ck(clk), .q(
        \pipeline/regfile/data[10][25] ) );
  dp_1 \pipeline/regfile/data_reg[10][26]  ( .ip(n9582), .ck(clk), .q(
        \pipeline/regfile/data[10][26] ) );
  dp_1 \pipeline/regfile/data_reg[10][27]  ( .ip(n9581), .ck(clk), .q(
        \pipeline/regfile/data[10][27] ) );
  dp_1 \pipeline/regfile/data_reg[10][28]  ( .ip(n9580), .ck(clk), .q(
        \pipeline/regfile/data[10][28] ) );
  dp_1 \pipeline/regfile/data_reg[10][29]  ( .ip(n9579), .ck(clk), .q(
        \pipeline/regfile/data[10][29] ) );
  dp_1 \pipeline/regfile/data_reg[10][30]  ( .ip(n9578), .ck(clk), .q(
        \pipeline/regfile/data[10][30] ) );
  dp_1 \pipeline/regfile/data_reg[10][31]  ( .ip(n9577), .ck(clk), .q(
        \pipeline/regfile/data[10][31] ) );
  dp_1 \pipeline/regfile/data_reg[11][0]  ( .ip(n9576), .ck(clk), .q(
        \pipeline/regfile/data[11][0] ) );
  dp_1 \pipeline/regfile/data_reg[11][1]  ( .ip(n9575), .ck(clk), .q(
        \pipeline/regfile/data[11][1] ) );
  dp_1 \pipeline/regfile/data_reg[11][2]  ( .ip(n9574), .ck(clk), .q(
        \pipeline/regfile/data[11][2] ) );
  dp_1 \pipeline/regfile/data_reg[11][3]  ( .ip(n9573), .ck(clk), .q(
        \pipeline/regfile/data[11][3] ) );
  dp_1 \pipeline/regfile/data_reg[11][4]  ( .ip(n9572), .ck(clk), .q(
        \pipeline/regfile/data[11][4] ) );
  dp_1 \pipeline/regfile/data_reg[11][5]  ( .ip(n9571), .ck(clk), .q(
        \pipeline/regfile/data[11][5] ) );
  dp_1 \pipeline/regfile/data_reg[11][6]  ( .ip(n9570), .ck(clk), .q(
        \pipeline/regfile/data[11][6] ) );
  dp_1 \pipeline/regfile/data_reg[11][7]  ( .ip(n9569), .ck(clk), .q(
        \pipeline/regfile/data[11][7] ) );
  dp_1 \pipeline/regfile/data_reg[11][8]  ( .ip(n9568), .ck(clk), .q(
        \pipeline/regfile/data[11][8] ) );
  dp_1 \pipeline/regfile/data_reg[11][9]  ( .ip(n9567), .ck(clk), .q(
        \pipeline/regfile/data[11][9] ) );
  dp_1 \pipeline/regfile/data_reg[11][10]  ( .ip(n9566), .ck(clk), .q(
        \pipeline/regfile/data[11][10] ) );
  dp_1 \pipeline/regfile/data_reg[11][11]  ( .ip(n9565), .ck(clk), .q(
        \pipeline/regfile/data[11][11] ) );
  dp_1 \pipeline/regfile/data_reg[11][12]  ( .ip(n9564), .ck(clk), .q(
        \pipeline/regfile/data[11][12] ) );
  dp_1 \pipeline/regfile/data_reg[11][13]  ( .ip(n9563), .ck(clk), .q(
        \pipeline/regfile/data[11][13] ) );
  dp_1 \pipeline/regfile/data_reg[11][14]  ( .ip(n9562), .ck(clk), .q(
        \pipeline/regfile/data[11][14] ) );
  dp_1 \pipeline/regfile/data_reg[11][15]  ( .ip(n9561), .ck(clk), .q(
        \pipeline/regfile/data[11][15] ) );
  dp_1 \pipeline/regfile/data_reg[11][16]  ( .ip(n9560), .ck(clk), .q(
        \pipeline/regfile/data[11][16] ) );
  dp_1 \pipeline/regfile/data_reg[11][17]  ( .ip(n9559), .ck(clk), .q(
        \pipeline/regfile/data[11][17] ) );
  dp_1 \pipeline/regfile/data_reg[11][18]  ( .ip(n9558), .ck(clk), .q(
        \pipeline/regfile/data[11][18] ) );
  dp_1 \pipeline/regfile/data_reg[11][19]  ( .ip(n9557), .ck(clk), .q(
        \pipeline/regfile/data[11][19] ) );
  dp_1 \pipeline/regfile/data_reg[11][20]  ( .ip(n9556), .ck(clk), .q(
        \pipeline/regfile/data[11][20] ) );
  dp_1 \pipeline/regfile/data_reg[11][21]  ( .ip(n9555), .ck(clk), .q(
        \pipeline/regfile/data[11][21] ) );
  dp_1 \pipeline/regfile/data_reg[11][22]  ( .ip(n9554), .ck(clk), .q(
        \pipeline/regfile/data[11][22] ) );
  dp_1 \pipeline/regfile/data_reg[11][23]  ( .ip(n9553), .ck(clk), .q(
        \pipeline/regfile/data[11][23] ) );
  dp_1 \pipeline/regfile/data_reg[11][24]  ( .ip(n9552), .ck(clk), .q(
        \pipeline/regfile/data[11][24] ) );
  dp_1 \pipeline/regfile/data_reg[11][25]  ( .ip(n9551), .ck(clk), .q(
        \pipeline/regfile/data[11][25] ) );
  dp_1 \pipeline/regfile/data_reg[11][26]  ( .ip(n9550), .ck(clk), .q(
        \pipeline/regfile/data[11][26] ) );
  dp_1 \pipeline/regfile/data_reg[11][27]  ( .ip(n9549), .ck(clk), .q(
        \pipeline/regfile/data[11][27] ) );
  dp_1 \pipeline/regfile/data_reg[11][28]  ( .ip(n9548), .ck(clk), .q(
        \pipeline/regfile/data[11][28] ) );
  dp_1 \pipeline/regfile/data_reg[11][29]  ( .ip(n9547), .ck(clk), .q(
        \pipeline/regfile/data[11][29] ) );
  dp_1 \pipeline/regfile/data_reg[11][30]  ( .ip(n9546), .ck(clk), .q(
        \pipeline/regfile/data[11][30] ) );
  dp_1 \pipeline/regfile/data_reg[11][31]  ( .ip(n9545), .ck(clk), .q(
        \pipeline/regfile/data[11][31] ) );
  dp_1 \pipeline/regfile/data_reg[12][0]  ( .ip(n9544), .ck(clk), .q(
        \pipeline/regfile/data[12][0] ) );
  dp_1 \pipeline/regfile/data_reg[12][1]  ( .ip(n9543), .ck(clk), .q(
        \pipeline/regfile/data[12][1] ) );
  dp_1 \pipeline/regfile/data_reg[12][2]  ( .ip(n9542), .ck(clk), .q(
        \pipeline/regfile/data[12][2] ) );
  dp_1 \pipeline/regfile/data_reg[12][3]  ( .ip(n9541), .ck(clk), .q(
        \pipeline/regfile/data[12][3] ) );
  dp_1 \pipeline/regfile/data_reg[12][4]  ( .ip(n9540), .ck(clk), .q(
        \pipeline/regfile/data[12][4] ) );
  dp_1 \pipeline/regfile/data_reg[12][5]  ( .ip(n9539), .ck(clk), .q(
        \pipeline/regfile/data[12][5] ) );
  dp_1 \pipeline/regfile/data_reg[12][6]  ( .ip(n9538), .ck(clk), .q(
        \pipeline/regfile/data[12][6] ) );
  dp_1 \pipeline/regfile/data_reg[12][7]  ( .ip(n9537), .ck(clk), .q(
        \pipeline/regfile/data[12][7] ) );
  dp_1 \pipeline/regfile/data_reg[12][8]  ( .ip(n9536), .ck(clk), .q(
        \pipeline/regfile/data[12][8] ) );
  dp_1 \pipeline/regfile/data_reg[12][9]  ( .ip(n9535), .ck(clk), .q(
        \pipeline/regfile/data[12][9] ) );
  dp_1 \pipeline/regfile/data_reg[12][10]  ( .ip(n9534), .ck(clk), .q(
        \pipeline/regfile/data[12][10] ) );
  dp_1 \pipeline/regfile/data_reg[12][11]  ( .ip(n9533), .ck(clk), .q(
        \pipeline/regfile/data[12][11] ) );
  dp_1 \pipeline/regfile/data_reg[12][12]  ( .ip(n9532), .ck(clk), .q(
        \pipeline/regfile/data[12][12] ) );
  dp_1 \pipeline/regfile/data_reg[12][13]  ( .ip(n9531), .ck(clk), .q(
        \pipeline/regfile/data[12][13] ) );
  dp_1 \pipeline/regfile/data_reg[12][14]  ( .ip(n9530), .ck(clk), .q(
        \pipeline/regfile/data[12][14] ) );
  dp_1 \pipeline/regfile/data_reg[12][15]  ( .ip(n9529), .ck(clk), .q(
        \pipeline/regfile/data[12][15] ) );
  dp_1 \pipeline/regfile/data_reg[12][16]  ( .ip(n9528), .ck(clk), .q(
        \pipeline/regfile/data[12][16] ) );
  dp_1 \pipeline/regfile/data_reg[12][17]  ( .ip(n9527), .ck(clk), .q(
        \pipeline/regfile/data[12][17] ) );
  dp_1 \pipeline/regfile/data_reg[12][18]  ( .ip(n9526), .ck(clk), .q(
        \pipeline/regfile/data[12][18] ) );
  dp_1 \pipeline/regfile/data_reg[12][19]  ( .ip(n9525), .ck(clk), .q(
        \pipeline/regfile/data[12][19] ) );
  dp_1 \pipeline/regfile/data_reg[12][20]  ( .ip(n9524), .ck(clk), .q(
        \pipeline/regfile/data[12][20] ) );
  dp_1 \pipeline/regfile/data_reg[12][21]  ( .ip(n9523), .ck(clk), .q(
        \pipeline/regfile/data[12][21] ) );
  dp_1 \pipeline/regfile/data_reg[12][22]  ( .ip(n9522), .ck(clk), .q(
        \pipeline/regfile/data[12][22] ) );
  dp_1 \pipeline/regfile/data_reg[12][23]  ( .ip(n9521), .ck(clk), .q(
        \pipeline/regfile/data[12][23] ) );
  dp_1 \pipeline/regfile/data_reg[12][24]  ( .ip(n9520), .ck(clk), .q(
        \pipeline/regfile/data[12][24] ) );
  dp_1 \pipeline/regfile/data_reg[12][25]  ( .ip(n9519), .ck(clk), .q(
        \pipeline/regfile/data[12][25] ) );
  dp_1 \pipeline/regfile/data_reg[12][26]  ( .ip(n9518), .ck(clk), .q(
        \pipeline/regfile/data[12][26] ) );
  dp_1 \pipeline/regfile/data_reg[12][27]  ( .ip(n9517), .ck(clk), .q(
        \pipeline/regfile/data[12][27] ) );
  dp_1 \pipeline/regfile/data_reg[12][28]  ( .ip(n9516), .ck(clk), .q(
        \pipeline/regfile/data[12][28] ) );
  dp_1 \pipeline/regfile/data_reg[12][29]  ( .ip(n9515), .ck(clk), .q(
        \pipeline/regfile/data[12][29] ) );
  dp_1 \pipeline/regfile/data_reg[12][30]  ( .ip(n9514), .ck(clk), .q(
        \pipeline/regfile/data[12][30] ) );
  dp_1 \pipeline/regfile/data_reg[12][31]  ( .ip(n9513), .ck(clk), .q(
        \pipeline/regfile/data[12][31] ) );
  dp_1 \pipeline/regfile/data_reg[13][0]  ( .ip(n9512), .ck(clk), .q(
        \pipeline/regfile/data[13][0] ) );
  dp_1 \pipeline/regfile/data_reg[13][1]  ( .ip(n9511), .ck(clk), .q(
        \pipeline/regfile/data[13][1] ) );
  dp_1 \pipeline/regfile/data_reg[13][2]  ( .ip(n9510), .ck(clk), .q(
        \pipeline/regfile/data[13][2] ) );
  dp_1 \pipeline/regfile/data_reg[13][3]  ( .ip(n9509), .ck(clk), .q(
        \pipeline/regfile/data[13][3] ) );
  dp_1 \pipeline/regfile/data_reg[13][4]  ( .ip(n9508), .ck(clk), .q(
        \pipeline/regfile/data[13][4] ) );
  dp_1 \pipeline/regfile/data_reg[13][5]  ( .ip(n9507), .ck(clk), .q(
        \pipeline/regfile/data[13][5] ) );
  dp_1 \pipeline/regfile/data_reg[13][6]  ( .ip(n9506), .ck(clk), .q(
        \pipeline/regfile/data[13][6] ) );
  dp_1 \pipeline/regfile/data_reg[13][7]  ( .ip(n9505), .ck(clk), .q(
        \pipeline/regfile/data[13][7] ) );
  dp_1 \pipeline/regfile/data_reg[13][8]  ( .ip(n9504), .ck(clk), .q(
        \pipeline/regfile/data[13][8] ) );
  dp_1 \pipeline/regfile/data_reg[13][9]  ( .ip(n9503), .ck(clk), .q(
        \pipeline/regfile/data[13][9] ) );
  dp_1 \pipeline/regfile/data_reg[13][10]  ( .ip(n9502), .ck(clk), .q(
        \pipeline/regfile/data[13][10] ) );
  dp_1 \pipeline/regfile/data_reg[13][11]  ( .ip(n9501), .ck(clk), .q(
        \pipeline/regfile/data[13][11] ) );
  dp_1 \pipeline/regfile/data_reg[13][12]  ( .ip(n9500), .ck(clk), .q(
        \pipeline/regfile/data[13][12] ) );
  dp_1 \pipeline/regfile/data_reg[13][13]  ( .ip(n9499), .ck(clk), .q(
        \pipeline/regfile/data[13][13] ) );
  dp_1 \pipeline/regfile/data_reg[13][14]  ( .ip(n9498), .ck(clk), .q(
        \pipeline/regfile/data[13][14] ) );
  dp_1 \pipeline/regfile/data_reg[13][15]  ( .ip(n9497), .ck(clk), .q(
        \pipeline/regfile/data[13][15] ) );
  dp_1 \pipeline/regfile/data_reg[13][16]  ( .ip(n9496), .ck(clk), .q(
        \pipeline/regfile/data[13][16] ) );
  dp_1 \pipeline/regfile/data_reg[13][17]  ( .ip(n9495), .ck(clk), .q(
        \pipeline/regfile/data[13][17] ) );
  dp_1 \pipeline/regfile/data_reg[13][18]  ( .ip(n9494), .ck(clk), .q(
        \pipeline/regfile/data[13][18] ) );
  dp_1 \pipeline/regfile/data_reg[13][19]  ( .ip(n9493), .ck(clk), .q(
        \pipeline/regfile/data[13][19] ) );
  dp_1 \pipeline/regfile/data_reg[13][20]  ( .ip(n9492), .ck(clk), .q(
        \pipeline/regfile/data[13][20] ) );
  dp_1 \pipeline/regfile/data_reg[13][21]  ( .ip(n9491), .ck(clk), .q(
        \pipeline/regfile/data[13][21] ) );
  dp_1 \pipeline/regfile/data_reg[13][22]  ( .ip(n9490), .ck(clk), .q(
        \pipeline/regfile/data[13][22] ) );
  dp_1 \pipeline/regfile/data_reg[13][23]  ( .ip(n9489), .ck(clk), .q(
        \pipeline/regfile/data[13][23] ) );
  dp_1 \pipeline/regfile/data_reg[13][24]  ( .ip(n9488), .ck(clk), .q(
        \pipeline/regfile/data[13][24] ) );
  dp_1 \pipeline/regfile/data_reg[13][25]  ( .ip(n9487), .ck(clk), .q(
        \pipeline/regfile/data[13][25] ) );
  dp_1 \pipeline/regfile/data_reg[13][26]  ( .ip(n9486), .ck(clk), .q(
        \pipeline/regfile/data[13][26] ) );
  dp_1 \pipeline/regfile/data_reg[13][27]  ( .ip(n9485), .ck(clk), .q(
        \pipeline/regfile/data[13][27] ) );
  dp_1 \pipeline/regfile/data_reg[13][28]  ( .ip(n9484), .ck(clk), .q(
        \pipeline/regfile/data[13][28] ) );
  dp_1 \pipeline/regfile/data_reg[13][29]  ( .ip(n9483), .ck(clk), .q(
        \pipeline/regfile/data[13][29] ) );
  dp_1 \pipeline/regfile/data_reg[13][30]  ( .ip(n9482), .ck(clk), .q(
        \pipeline/regfile/data[13][30] ) );
  dp_1 \pipeline/regfile/data_reg[13][31]  ( .ip(n9481), .ck(clk), .q(
        \pipeline/regfile/data[13][31] ) );
  dp_1 \pipeline/regfile/data_reg[14][0]  ( .ip(n9480), .ck(clk), .q(
        \pipeline/regfile/data[14][0] ) );
  dp_1 \pipeline/regfile/data_reg[14][1]  ( .ip(n9479), .ck(clk), .q(
        \pipeline/regfile/data[14][1] ) );
  dp_1 \pipeline/regfile/data_reg[14][2]  ( .ip(n9478), .ck(clk), .q(
        \pipeline/regfile/data[14][2] ) );
  dp_1 \pipeline/regfile/data_reg[14][3]  ( .ip(n9477), .ck(clk), .q(
        \pipeline/regfile/data[14][3] ) );
  dp_1 \pipeline/regfile/data_reg[14][4]  ( .ip(n9476), .ck(clk), .q(
        \pipeline/regfile/data[14][4] ) );
  dp_1 \pipeline/regfile/data_reg[14][5]  ( .ip(n9475), .ck(clk), .q(
        \pipeline/regfile/data[14][5] ) );
  dp_1 \pipeline/regfile/data_reg[14][6]  ( .ip(n9474), .ck(clk), .q(
        \pipeline/regfile/data[14][6] ) );
  dp_1 \pipeline/regfile/data_reg[14][7]  ( .ip(n9473), .ck(clk), .q(
        \pipeline/regfile/data[14][7] ) );
  dp_1 \pipeline/regfile/data_reg[14][8]  ( .ip(n9472), .ck(clk), .q(
        \pipeline/regfile/data[14][8] ) );
  dp_1 \pipeline/regfile/data_reg[14][9]  ( .ip(n9471), .ck(clk), .q(
        \pipeline/regfile/data[14][9] ) );
  dp_1 \pipeline/regfile/data_reg[14][10]  ( .ip(n9470), .ck(clk), .q(
        \pipeline/regfile/data[14][10] ) );
  dp_1 \pipeline/regfile/data_reg[14][11]  ( .ip(n9469), .ck(clk), .q(
        \pipeline/regfile/data[14][11] ) );
  dp_1 \pipeline/regfile/data_reg[14][12]  ( .ip(n9468), .ck(clk), .q(
        \pipeline/regfile/data[14][12] ) );
  dp_1 \pipeline/regfile/data_reg[14][13]  ( .ip(n9467), .ck(clk), .q(
        \pipeline/regfile/data[14][13] ) );
  dp_1 \pipeline/regfile/data_reg[14][14]  ( .ip(n9466), .ck(clk), .q(
        \pipeline/regfile/data[14][14] ) );
  dp_1 \pipeline/regfile/data_reg[14][15]  ( .ip(n9465), .ck(clk), .q(
        \pipeline/regfile/data[14][15] ) );
  dp_1 \pipeline/regfile/data_reg[14][16]  ( .ip(n9464), .ck(clk), .q(
        \pipeline/regfile/data[14][16] ) );
  dp_1 \pipeline/regfile/data_reg[14][17]  ( .ip(n9463), .ck(clk), .q(
        \pipeline/regfile/data[14][17] ) );
  dp_1 \pipeline/regfile/data_reg[14][18]  ( .ip(n9462), .ck(clk), .q(
        \pipeline/regfile/data[14][18] ) );
  dp_1 \pipeline/regfile/data_reg[14][19]  ( .ip(n9461), .ck(clk), .q(
        \pipeline/regfile/data[14][19] ) );
  dp_1 \pipeline/regfile/data_reg[14][20]  ( .ip(n9460), .ck(clk), .q(
        \pipeline/regfile/data[14][20] ) );
  dp_1 \pipeline/regfile/data_reg[14][21]  ( .ip(n9459), .ck(clk), .q(
        \pipeline/regfile/data[14][21] ) );
  dp_1 \pipeline/regfile/data_reg[14][22]  ( .ip(n9458), .ck(clk), .q(
        \pipeline/regfile/data[14][22] ) );
  dp_1 \pipeline/regfile/data_reg[14][23]  ( .ip(n9457), .ck(clk), .q(
        \pipeline/regfile/data[14][23] ) );
  dp_1 \pipeline/regfile/data_reg[14][24]  ( .ip(n9456), .ck(clk), .q(
        \pipeline/regfile/data[14][24] ) );
  dp_1 \pipeline/regfile/data_reg[14][25]  ( .ip(n9455), .ck(clk), .q(
        \pipeline/regfile/data[14][25] ) );
  dp_1 \pipeline/regfile/data_reg[14][26]  ( .ip(n9454), .ck(clk), .q(
        \pipeline/regfile/data[14][26] ) );
  dp_1 \pipeline/regfile/data_reg[14][27]  ( .ip(n9453), .ck(clk), .q(
        \pipeline/regfile/data[14][27] ) );
  dp_1 \pipeline/regfile/data_reg[14][28]  ( .ip(n9452), .ck(clk), .q(
        \pipeline/regfile/data[14][28] ) );
  dp_1 \pipeline/regfile/data_reg[14][29]  ( .ip(n9451), .ck(clk), .q(
        \pipeline/regfile/data[14][29] ) );
  dp_1 \pipeline/regfile/data_reg[14][30]  ( .ip(n9450), .ck(clk), .q(
        \pipeline/regfile/data[14][30] ) );
  dp_1 \pipeline/regfile/data_reg[14][31]  ( .ip(n9449), .ck(clk), .q(
        \pipeline/regfile/data[14][31] ) );
  dp_1 \pipeline/regfile/data_reg[15][0]  ( .ip(n9448), .ck(clk), .q(
        \pipeline/regfile/data[15][0] ) );
  dp_1 \pipeline/regfile/data_reg[15][1]  ( .ip(n9447), .ck(clk), .q(
        \pipeline/regfile/data[15][1] ) );
  dp_1 \pipeline/regfile/data_reg[15][2]  ( .ip(n9446), .ck(clk), .q(
        \pipeline/regfile/data[15][2] ) );
  dp_1 \pipeline/regfile/data_reg[15][3]  ( .ip(n9445), .ck(clk), .q(
        \pipeline/regfile/data[15][3] ) );
  dp_1 \pipeline/regfile/data_reg[15][4]  ( .ip(n9444), .ck(clk), .q(
        \pipeline/regfile/data[15][4] ) );
  dp_1 \pipeline/regfile/data_reg[15][5]  ( .ip(n9443), .ck(clk), .q(
        \pipeline/regfile/data[15][5] ) );
  dp_1 \pipeline/regfile/data_reg[15][6]  ( .ip(n9442), .ck(clk), .q(
        \pipeline/regfile/data[15][6] ) );
  dp_1 \pipeline/regfile/data_reg[15][7]  ( .ip(n9441), .ck(clk), .q(
        \pipeline/regfile/data[15][7] ) );
  dp_1 \pipeline/regfile/data_reg[15][8]  ( .ip(n9440), .ck(clk), .q(
        \pipeline/regfile/data[15][8] ) );
  dp_1 \pipeline/regfile/data_reg[15][9]  ( .ip(n9439), .ck(clk), .q(
        \pipeline/regfile/data[15][9] ) );
  dp_1 \pipeline/regfile/data_reg[15][10]  ( .ip(n9438), .ck(clk), .q(
        \pipeline/regfile/data[15][10] ) );
  dp_1 \pipeline/regfile/data_reg[15][11]  ( .ip(n9437), .ck(clk), .q(
        \pipeline/regfile/data[15][11] ) );
  dp_1 \pipeline/regfile/data_reg[15][12]  ( .ip(n9436), .ck(clk), .q(
        \pipeline/regfile/data[15][12] ) );
  dp_1 \pipeline/regfile/data_reg[15][13]  ( .ip(n9435), .ck(clk), .q(
        \pipeline/regfile/data[15][13] ) );
  dp_1 \pipeline/regfile/data_reg[15][14]  ( .ip(n9434), .ck(clk), .q(
        \pipeline/regfile/data[15][14] ) );
  dp_1 \pipeline/regfile/data_reg[15][15]  ( .ip(n9433), .ck(clk), .q(
        \pipeline/regfile/data[15][15] ) );
  dp_1 \pipeline/regfile/data_reg[15][16]  ( .ip(n9432), .ck(clk), .q(
        \pipeline/regfile/data[15][16] ) );
  dp_1 \pipeline/regfile/data_reg[15][17]  ( .ip(n9431), .ck(clk), .q(
        \pipeline/regfile/data[15][17] ) );
  dp_1 \pipeline/regfile/data_reg[15][18]  ( .ip(n9430), .ck(clk), .q(
        \pipeline/regfile/data[15][18] ) );
  dp_1 \pipeline/regfile/data_reg[15][19]  ( .ip(n9429), .ck(clk), .q(
        \pipeline/regfile/data[15][19] ) );
  dp_1 \pipeline/regfile/data_reg[15][20]  ( .ip(n9428), .ck(clk), .q(
        \pipeline/regfile/data[15][20] ) );
  dp_1 \pipeline/regfile/data_reg[15][21]  ( .ip(n9427), .ck(clk), .q(
        \pipeline/regfile/data[15][21] ) );
  dp_1 \pipeline/regfile/data_reg[15][22]  ( .ip(n9426), .ck(clk), .q(
        \pipeline/regfile/data[15][22] ) );
  dp_1 \pipeline/regfile/data_reg[15][23]  ( .ip(n9425), .ck(clk), .q(
        \pipeline/regfile/data[15][23] ) );
  dp_1 \pipeline/regfile/data_reg[15][24]  ( .ip(n9424), .ck(clk), .q(
        \pipeline/regfile/data[15][24] ) );
  dp_1 \pipeline/regfile/data_reg[15][25]  ( .ip(n9423), .ck(clk), .q(
        \pipeline/regfile/data[15][25] ) );
  dp_1 \pipeline/regfile/data_reg[15][26]  ( .ip(n9422), .ck(clk), .q(
        \pipeline/regfile/data[15][26] ) );
  dp_1 \pipeline/regfile/data_reg[15][27]  ( .ip(n9421), .ck(clk), .q(
        \pipeline/regfile/data[15][27] ) );
  dp_1 \pipeline/regfile/data_reg[15][28]  ( .ip(n9420), .ck(clk), .q(
        \pipeline/regfile/data[15][28] ) );
  dp_1 \pipeline/regfile/data_reg[15][29]  ( .ip(n9419), .ck(clk), .q(
        \pipeline/regfile/data[15][29] ) );
  dp_1 \pipeline/regfile/data_reg[15][30]  ( .ip(n9418), .ck(clk), .q(
        \pipeline/regfile/data[15][30] ) );
  dp_1 \pipeline/regfile/data_reg[15][31]  ( .ip(n9417), .ck(clk), .q(
        \pipeline/regfile/data[15][31] ) );
  dp_1 \pipeline/regfile/data_reg[16][0]  ( .ip(n9416), .ck(clk), .q(
        \pipeline/regfile/data[16][0] ) );
  dp_1 \pipeline/regfile/data_reg[16][1]  ( .ip(n9415), .ck(clk), .q(
        \pipeline/regfile/data[16][1] ) );
  dp_1 \pipeline/regfile/data_reg[16][2]  ( .ip(n9414), .ck(clk), .q(
        \pipeline/regfile/data[16][2] ) );
  dp_1 \pipeline/regfile/data_reg[16][3]  ( .ip(n9413), .ck(clk), .q(
        \pipeline/regfile/data[16][3] ) );
  dp_1 \pipeline/regfile/data_reg[16][4]  ( .ip(n9412), .ck(clk), .q(
        \pipeline/regfile/data[16][4] ) );
  dp_1 \pipeline/regfile/data_reg[16][5]  ( .ip(n9411), .ck(clk), .q(
        \pipeline/regfile/data[16][5] ) );
  dp_1 \pipeline/regfile/data_reg[16][6]  ( .ip(n9410), .ck(clk), .q(
        \pipeline/regfile/data[16][6] ) );
  dp_1 \pipeline/regfile/data_reg[16][7]  ( .ip(n9409), .ck(clk), .q(
        \pipeline/regfile/data[16][7] ) );
  dp_1 \pipeline/regfile/data_reg[16][8]  ( .ip(n9408), .ck(clk), .q(
        \pipeline/regfile/data[16][8] ) );
  dp_1 \pipeline/regfile/data_reg[16][9]  ( .ip(n9407), .ck(clk), .q(
        \pipeline/regfile/data[16][9] ) );
  dp_1 \pipeline/regfile/data_reg[16][10]  ( .ip(n9406), .ck(clk), .q(
        \pipeline/regfile/data[16][10] ) );
  dp_1 \pipeline/regfile/data_reg[16][11]  ( .ip(n9405), .ck(clk), .q(
        \pipeline/regfile/data[16][11] ) );
  dp_1 \pipeline/regfile/data_reg[16][12]  ( .ip(n9404), .ck(clk), .q(
        \pipeline/regfile/data[16][12] ) );
  dp_1 \pipeline/regfile/data_reg[16][13]  ( .ip(n9403), .ck(clk), .q(
        \pipeline/regfile/data[16][13] ) );
  dp_1 \pipeline/regfile/data_reg[16][14]  ( .ip(n9402), .ck(clk), .q(
        \pipeline/regfile/data[16][14] ) );
  dp_1 \pipeline/regfile/data_reg[16][15]  ( .ip(n9401), .ck(clk), .q(
        \pipeline/regfile/data[16][15] ) );
  dp_1 \pipeline/regfile/data_reg[16][16]  ( .ip(n9400), .ck(clk), .q(
        \pipeline/regfile/data[16][16] ) );
  dp_1 \pipeline/regfile/data_reg[16][17]  ( .ip(n9399), .ck(clk), .q(
        \pipeline/regfile/data[16][17] ) );
  dp_1 \pipeline/regfile/data_reg[16][18]  ( .ip(n9398), .ck(clk), .q(
        \pipeline/regfile/data[16][18] ) );
  dp_1 \pipeline/regfile/data_reg[16][19]  ( .ip(n9397), .ck(clk), .q(
        \pipeline/regfile/data[16][19] ) );
  dp_1 \pipeline/regfile/data_reg[16][20]  ( .ip(n9396), .ck(clk), .q(
        \pipeline/regfile/data[16][20] ) );
  dp_1 \pipeline/regfile/data_reg[16][21]  ( .ip(n9395), .ck(clk), .q(
        \pipeline/regfile/data[16][21] ) );
  dp_1 \pipeline/regfile/data_reg[16][22]  ( .ip(n9394), .ck(clk), .q(
        \pipeline/regfile/data[16][22] ) );
  dp_1 \pipeline/regfile/data_reg[16][23]  ( .ip(n9393), .ck(clk), .q(
        \pipeline/regfile/data[16][23] ) );
  dp_1 \pipeline/regfile/data_reg[16][24]  ( .ip(n9392), .ck(clk), .q(
        \pipeline/regfile/data[16][24] ) );
  dp_1 \pipeline/regfile/data_reg[16][25]  ( .ip(n9391), .ck(clk), .q(
        \pipeline/regfile/data[16][25] ) );
  dp_1 \pipeline/regfile/data_reg[16][26]  ( .ip(n9390), .ck(clk), .q(
        \pipeline/regfile/data[16][26] ) );
  dp_1 \pipeline/regfile/data_reg[16][27]  ( .ip(n9389), .ck(clk), .q(
        \pipeline/regfile/data[16][27] ) );
  dp_1 \pipeline/regfile/data_reg[16][28]  ( .ip(n9388), .ck(clk), .q(
        \pipeline/regfile/data[16][28] ) );
  dp_1 \pipeline/regfile/data_reg[16][29]  ( .ip(n9387), .ck(clk), .q(
        \pipeline/regfile/data[16][29] ) );
  dp_1 \pipeline/regfile/data_reg[16][30]  ( .ip(n9386), .ck(clk), .q(
        \pipeline/regfile/data[16][30] ) );
  dp_1 \pipeline/regfile/data_reg[16][31]  ( .ip(n9385), .ck(clk), .q(
        \pipeline/regfile/data[16][31] ) );
  dp_1 \pipeline/regfile/data_reg[17][0]  ( .ip(n9384), .ck(clk), .q(
        \pipeline/regfile/data[17][0] ) );
  dp_1 \pipeline/regfile/data_reg[17][1]  ( .ip(n9383), .ck(clk), .q(
        \pipeline/regfile/data[17][1] ) );
  dp_1 \pipeline/regfile/data_reg[17][2]  ( .ip(n9382), .ck(clk), .q(
        \pipeline/regfile/data[17][2] ) );
  dp_1 \pipeline/regfile/data_reg[17][3]  ( .ip(n9381), .ck(clk), .q(
        \pipeline/regfile/data[17][3] ) );
  dp_1 \pipeline/regfile/data_reg[17][4]  ( .ip(n9380), .ck(clk), .q(
        \pipeline/regfile/data[17][4] ) );
  dp_1 \pipeline/regfile/data_reg[17][5]  ( .ip(n9379), .ck(clk), .q(
        \pipeline/regfile/data[17][5] ) );
  dp_1 \pipeline/regfile/data_reg[17][6]  ( .ip(n9378), .ck(clk), .q(
        \pipeline/regfile/data[17][6] ) );
  dp_1 \pipeline/regfile/data_reg[17][7]  ( .ip(n9377), .ck(clk), .q(
        \pipeline/regfile/data[17][7] ) );
  dp_1 \pipeline/regfile/data_reg[17][8]  ( .ip(n9376), .ck(clk), .q(
        \pipeline/regfile/data[17][8] ) );
  dp_1 \pipeline/regfile/data_reg[17][9]  ( .ip(n9375), .ck(clk), .q(
        \pipeline/regfile/data[17][9] ) );
  dp_1 \pipeline/regfile/data_reg[17][10]  ( .ip(n9374), .ck(clk), .q(
        \pipeline/regfile/data[17][10] ) );
  dp_1 \pipeline/regfile/data_reg[17][11]  ( .ip(n9373), .ck(clk), .q(
        \pipeline/regfile/data[17][11] ) );
  dp_1 \pipeline/regfile/data_reg[17][12]  ( .ip(n9372), .ck(clk), .q(
        \pipeline/regfile/data[17][12] ) );
  dp_1 \pipeline/regfile/data_reg[17][13]  ( .ip(n9371), .ck(clk), .q(
        \pipeline/regfile/data[17][13] ) );
  dp_1 \pipeline/regfile/data_reg[17][14]  ( .ip(n9370), .ck(clk), .q(
        \pipeline/regfile/data[17][14] ) );
  dp_1 \pipeline/regfile/data_reg[17][15]  ( .ip(n9369), .ck(clk), .q(
        \pipeline/regfile/data[17][15] ) );
  dp_1 \pipeline/regfile/data_reg[17][16]  ( .ip(n9368), .ck(clk), .q(
        \pipeline/regfile/data[17][16] ) );
  dp_1 \pipeline/regfile/data_reg[17][17]  ( .ip(n9367), .ck(clk), .q(
        \pipeline/regfile/data[17][17] ) );
  dp_1 \pipeline/regfile/data_reg[17][18]  ( .ip(n9366), .ck(clk), .q(
        \pipeline/regfile/data[17][18] ) );
  dp_1 \pipeline/regfile/data_reg[17][19]  ( .ip(n9365), .ck(clk), .q(
        \pipeline/regfile/data[17][19] ) );
  dp_1 \pipeline/regfile/data_reg[17][20]  ( .ip(n9364), .ck(clk), .q(
        \pipeline/regfile/data[17][20] ) );
  dp_1 \pipeline/regfile/data_reg[17][21]  ( .ip(n9363), .ck(clk), .q(
        \pipeline/regfile/data[17][21] ) );
  dp_1 \pipeline/regfile/data_reg[17][22]  ( .ip(n9362), .ck(clk), .q(
        \pipeline/regfile/data[17][22] ) );
  dp_1 \pipeline/regfile/data_reg[17][23]  ( .ip(n9361), .ck(clk), .q(
        \pipeline/regfile/data[17][23] ) );
  dp_1 \pipeline/regfile/data_reg[17][24]  ( .ip(n9360), .ck(clk), .q(
        \pipeline/regfile/data[17][24] ) );
  dp_1 \pipeline/regfile/data_reg[17][25]  ( .ip(n9359), .ck(clk), .q(
        \pipeline/regfile/data[17][25] ) );
  dp_1 \pipeline/regfile/data_reg[17][26]  ( .ip(n9358), .ck(clk), .q(
        \pipeline/regfile/data[17][26] ) );
  dp_1 \pipeline/regfile/data_reg[17][27]  ( .ip(n9357), .ck(clk), .q(
        \pipeline/regfile/data[17][27] ) );
  dp_1 \pipeline/regfile/data_reg[17][28]  ( .ip(n9356), .ck(clk), .q(
        \pipeline/regfile/data[17][28] ) );
  dp_1 \pipeline/regfile/data_reg[17][29]  ( .ip(n9355), .ck(clk), .q(
        \pipeline/regfile/data[17][29] ) );
  dp_1 \pipeline/regfile/data_reg[17][30]  ( .ip(n9354), .ck(clk), .q(
        \pipeline/regfile/data[17][30] ) );
  dp_1 \pipeline/regfile/data_reg[17][31]  ( .ip(n9353), .ck(clk), .q(
        \pipeline/regfile/data[17][31] ) );
  dp_1 \pipeline/regfile/data_reg[18][0]  ( .ip(n9352), .ck(clk), .q(
        \pipeline/regfile/data[18][0] ) );
  dp_1 \pipeline/regfile/data_reg[18][1]  ( .ip(n9351), .ck(clk), .q(
        \pipeline/regfile/data[18][1] ) );
  dp_1 \pipeline/regfile/data_reg[18][2]  ( .ip(n9350), .ck(clk), .q(
        \pipeline/regfile/data[18][2] ) );
  dp_1 \pipeline/regfile/data_reg[18][3]  ( .ip(n9349), .ck(clk), .q(
        \pipeline/regfile/data[18][3] ) );
  dp_1 \pipeline/regfile/data_reg[18][4]  ( .ip(n9348), .ck(clk), .q(
        \pipeline/regfile/data[18][4] ) );
  dp_1 \pipeline/regfile/data_reg[18][5]  ( .ip(n9347), .ck(clk), .q(
        \pipeline/regfile/data[18][5] ) );
  dp_1 \pipeline/regfile/data_reg[18][6]  ( .ip(n9346), .ck(clk), .q(
        \pipeline/regfile/data[18][6] ) );
  dp_1 \pipeline/regfile/data_reg[18][7]  ( .ip(n9345), .ck(clk), .q(
        \pipeline/regfile/data[18][7] ) );
  dp_1 \pipeline/regfile/data_reg[18][8]  ( .ip(n9344), .ck(clk), .q(
        \pipeline/regfile/data[18][8] ) );
  dp_1 \pipeline/regfile/data_reg[18][9]  ( .ip(n9343), .ck(clk), .q(
        \pipeline/regfile/data[18][9] ) );
  dp_1 \pipeline/regfile/data_reg[18][10]  ( .ip(n9342), .ck(clk), .q(
        \pipeline/regfile/data[18][10] ) );
  dp_1 \pipeline/regfile/data_reg[18][11]  ( .ip(n9341), .ck(clk), .q(
        \pipeline/regfile/data[18][11] ) );
  dp_1 \pipeline/regfile/data_reg[18][12]  ( .ip(n9340), .ck(clk), .q(
        \pipeline/regfile/data[18][12] ) );
  dp_1 \pipeline/regfile/data_reg[18][13]  ( .ip(n9339), .ck(clk), .q(
        \pipeline/regfile/data[18][13] ) );
  dp_1 \pipeline/regfile/data_reg[18][14]  ( .ip(n9338), .ck(clk), .q(
        \pipeline/regfile/data[18][14] ) );
  dp_1 \pipeline/regfile/data_reg[18][15]  ( .ip(n9337), .ck(clk), .q(
        \pipeline/regfile/data[18][15] ) );
  dp_1 \pipeline/regfile/data_reg[18][16]  ( .ip(n9336), .ck(clk), .q(
        \pipeline/regfile/data[18][16] ) );
  dp_1 \pipeline/regfile/data_reg[18][17]  ( .ip(n9335), .ck(clk), .q(
        \pipeline/regfile/data[18][17] ) );
  dp_1 \pipeline/regfile/data_reg[18][18]  ( .ip(n9334), .ck(clk), .q(
        \pipeline/regfile/data[18][18] ) );
  dp_1 \pipeline/regfile/data_reg[18][19]  ( .ip(n9333), .ck(clk), .q(
        \pipeline/regfile/data[18][19] ) );
  dp_1 \pipeline/regfile/data_reg[18][20]  ( .ip(n9332), .ck(clk), .q(
        \pipeline/regfile/data[18][20] ) );
  dp_1 \pipeline/regfile/data_reg[18][21]  ( .ip(n9331), .ck(clk), .q(
        \pipeline/regfile/data[18][21] ) );
  dp_1 \pipeline/regfile/data_reg[18][22]  ( .ip(n9330), .ck(clk), .q(
        \pipeline/regfile/data[18][22] ) );
  dp_1 \pipeline/regfile/data_reg[18][23]  ( .ip(n9329), .ck(clk), .q(
        \pipeline/regfile/data[18][23] ) );
  dp_1 \pipeline/regfile/data_reg[18][24]  ( .ip(n9328), .ck(clk), .q(
        \pipeline/regfile/data[18][24] ) );
  dp_1 \pipeline/regfile/data_reg[18][25]  ( .ip(n9327), .ck(clk), .q(
        \pipeline/regfile/data[18][25] ) );
  dp_1 \pipeline/regfile/data_reg[18][26]  ( .ip(n9326), .ck(clk), .q(
        \pipeline/regfile/data[18][26] ) );
  dp_1 \pipeline/regfile/data_reg[18][27]  ( .ip(n9325), .ck(clk), .q(
        \pipeline/regfile/data[18][27] ) );
  dp_1 \pipeline/regfile/data_reg[18][28]  ( .ip(n9324), .ck(clk), .q(
        \pipeline/regfile/data[18][28] ) );
  dp_1 \pipeline/regfile/data_reg[18][29]  ( .ip(n9323), .ck(clk), .q(
        \pipeline/regfile/data[18][29] ) );
  dp_1 \pipeline/regfile/data_reg[18][30]  ( .ip(n9322), .ck(clk), .q(
        \pipeline/regfile/data[18][30] ) );
  dp_1 \pipeline/regfile/data_reg[18][31]  ( .ip(n9321), .ck(clk), .q(
        \pipeline/regfile/data[18][31] ) );
  dp_1 \pipeline/regfile/data_reg[19][0]  ( .ip(n9320), .ck(clk), .q(
        \pipeline/regfile/data[19][0] ) );
  dp_1 \pipeline/regfile/data_reg[19][1]  ( .ip(n9319), .ck(clk), .q(
        \pipeline/regfile/data[19][1] ) );
  dp_1 \pipeline/regfile/data_reg[19][2]  ( .ip(n9318), .ck(clk), .q(
        \pipeline/regfile/data[19][2] ) );
  dp_1 \pipeline/regfile/data_reg[19][3]  ( .ip(n9317), .ck(clk), .q(
        \pipeline/regfile/data[19][3] ) );
  dp_1 \pipeline/regfile/data_reg[19][4]  ( .ip(n9316), .ck(clk), .q(
        \pipeline/regfile/data[19][4] ) );
  dp_1 \pipeline/regfile/data_reg[19][5]  ( .ip(n9315), .ck(clk), .q(
        \pipeline/regfile/data[19][5] ) );
  dp_1 \pipeline/regfile/data_reg[19][6]  ( .ip(n9314), .ck(clk), .q(
        \pipeline/regfile/data[19][6] ) );
  dp_1 \pipeline/regfile/data_reg[19][7]  ( .ip(n9313), .ck(clk), .q(
        \pipeline/regfile/data[19][7] ) );
  dp_1 \pipeline/regfile/data_reg[19][8]  ( .ip(n9312), .ck(clk), .q(
        \pipeline/regfile/data[19][8] ) );
  dp_1 \pipeline/regfile/data_reg[19][9]  ( .ip(n9311), .ck(clk), .q(
        \pipeline/regfile/data[19][9] ) );
  dp_1 \pipeline/regfile/data_reg[19][10]  ( .ip(n9310), .ck(clk), .q(
        \pipeline/regfile/data[19][10] ) );
  dp_1 \pipeline/regfile/data_reg[19][11]  ( .ip(n9309), .ck(clk), .q(
        \pipeline/regfile/data[19][11] ) );
  dp_1 \pipeline/regfile/data_reg[19][12]  ( .ip(n9308), .ck(clk), .q(
        \pipeline/regfile/data[19][12] ) );
  dp_1 \pipeline/regfile/data_reg[19][13]  ( .ip(n9307), .ck(clk), .q(
        \pipeline/regfile/data[19][13] ) );
  dp_1 \pipeline/regfile/data_reg[19][14]  ( .ip(n9306), .ck(clk), .q(
        \pipeline/regfile/data[19][14] ) );
  dp_1 \pipeline/regfile/data_reg[19][15]  ( .ip(n9305), .ck(clk), .q(
        \pipeline/regfile/data[19][15] ) );
  dp_1 \pipeline/regfile/data_reg[19][16]  ( .ip(n9304), .ck(clk), .q(
        \pipeline/regfile/data[19][16] ) );
  dp_1 \pipeline/regfile/data_reg[19][17]  ( .ip(n9303), .ck(clk), .q(
        \pipeline/regfile/data[19][17] ) );
  dp_1 \pipeline/regfile/data_reg[19][18]  ( .ip(n9302), .ck(clk), .q(
        \pipeline/regfile/data[19][18] ) );
  dp_1 \pipeline/regfile/data_reg[19][19]  ( .ip(n9301), .ck(clk), .q(
        \pipeline/regfile/data[19][19] ) );
  dp_1 \pipeline/regfile/data_reg[19][20]  ( .ip(n9300), .ck(clk), .q(
        \pipeline/regfile/data[19][20] ) );
  dp_1 \pipeline/regfile/data_reg[19][21]  ( .ip(n9299), .ck(clk), .q(
        \pipeline/regfile/data[19][21] ) );
  dp_1 \pipeline/regfile/data_reg[19][22]  ( .ip(n9298), .ck(clk), .q(
        \pipeline/regfile/data[19][22] ) );
  dp_1 \pipeline/regfile/data_reg[19][23]  ( .ip(n9297), .ck(clk), .q(
        \pipeline/regfile/data[19][23] ) );
  dp_1 \pipeline/regfile/data_reg[19][24]  ( .ip(n9296), .ck(clk), .q(
        \pipeline/regfile/data[19][24] ) );
  dp_1 \pipeline/regfile/data_reg[19][25]  ( .ip(n9295), .ck(clk), .q(
        \pipeline/regfile/data[19][25] ) );
  dp_1 \pipeline/regfile/data_reg[19][26]  ( .ip(n9294), .ck(clk), .q(
        \pipeline/regfile/data[19][26] ) );
  dp_1 \pipeline/regfile/data_reg[19][27]  ( .ip(n9293), .ck(clk), .q(
        \pipeline/regfile/data[19][27] ) );
  dp_1 \pipeline/regfile/data_reg[19][28]  ( .ip(n9292), .ck(clk), .q(
        \pipeline/regfile/data[19][28] ) );
  dp_1 \pipeline/regfile/data_reg[19][29]  ( .ip(n9291), .ck(clk), .q(
        \pipeline/regfile/data[19][29] ) );
  dp_1 \pipeline/regfile/data_reg[19][30]  ( .ip(n9290), .ck(clk), .q(
        \pipeline/regfile/data[19][30] ) );
  dp_1 \pipeline/regfile/data_reg[19][31]  ( .ip(n9289), .ck(clk), .q(
        \pipeline/regfile/data[19][31] ) );
  dp_1 \pipeline/regfile/data_reg[20][0]  ( .ip(n9288), .ck(clk), .q(
        \pipeline/regfile/data[20][0] ) );
  dp_1 \pipeline/regfile/data_reg[20][1]  ( .ip(n9287), .ck(clk), .q(
        \pipeline/regfile/data[20][1] ) );
  dp_1 \pipeline/regfile/data_reg[20][2]  ( .ip(n9286), .ck(clk), .q(
        \pipeline/regfile/data[20][2] ) );
  dp_1 \pipeline/regfile/data_reg[20][3]  ( .ip(n9285), .ck(clk), .q(
        \pipeline/regfile/data[20][3] ) );
  dp_1 \pipeline/regfile/data_reg[20][4]  ( .ip(n9284), .ck(clk), .q(
        \pipeline/regfile/data[20][4] ) );
  dp_1 \pipeline/regfile/data_reg[20][5]  ( .ip(n9283), .ck(clk), .q(
        \pipeline/regfile/data[20][5] ) );
  dp_1 \pipeline/regfile/data_reg[20][6]  ( .ip(n9282), .ck(clk), .q(
        \pipeline/regfile/data[20][6] ) );
  dp_1 \pipeline/regfile/data_reg[20][7]  ( .ip(n9281), .ck(clk), .q(
        \pipeline/regfile/data[20][7] ) );
  dp_1 \pipeline/regfile/data_reg[20][8]  ( .ip(n9280), .ck(clk), .q(
        \pipeline/regfile/data[20][8] ) );
  dp_1 \pipeline/regfile/data_reg[20][9]  ( .ip(n9279), .ck(clk), .q(
        \pipeline/regfile/data[20][9] ) );
  dp_1 \pipeline/regfile/data_reg[20][10]  ( .ip(n9278), .ck(clk), .q(
        \pipeline/regfile/data[20][10] ) );
  dp_1 \pipeline/regfile/data_reg[20][11]  ( .ip(n9277), .ck(clk), .q(
        \pipeline/regfile/data[20][11] ) );
  dp_1 \pipeline/regfile/data_reg[20][12]  ( .ip(n9276), .ck(clk), .q(
        \pipeline/regfile/data[20][12] ) );
  dp_1 \pipeline/regfile/data_reg[20][13]  ( .ip(n9275), .ck(clk), .q(
        \pipeline/regfile/data[20][13] ) );
  dp_1 \pipeline/regfile/data_reg[20][14]  ( .ip(n9274), .ck(clk), .q(
        \pipeline/regfile/data[20][14] ) );
  dp_1 \pipeline/regfile/data_reg[20][15]  ( .ip(n9273), .ck(clk), .q(
        \pipeline/regfile/data[20][15] ) );
  dp_1 \pipeline/regfile/data_reg[20][16]  ( .ip(n9272), .ck(clk), .q(
        \pipeline/regfile/data[20][16] ) );
  dp_1 \pipeline/regfile/data_reg[20][17]  ( .ip(n9271), .ck(clk), .q(
        \pipeline/regfile/data[20][17] ) );
  dp_1 \pipeline/regfile/data_reg[20][18]  ( .ip(n9270), .ck(clk), .q(
        \pipeline/regfile/data[20][18] ) );
  dp_1 \pipeline/regfile/data_reg[20][19]  ( .ip(n9269), .ck(clk), .q(
        \pipeline/regfile/data[20][19] ) );
  dp_1 \pipeline/regfile/data_reg[20][20]  ( .ip(n9268), .ck(clk), .q(
        \pipeline/regfile/data[20][20] ) );
  dp_1 \pipeline/regfile/data_reg[20][21]  ( .ip(n9267), .ck(clk), .q(
        \pipeline/regfile/data[20][21] ) );
  dp_1 \pipeline/regfile/data_reg[20][22]  ( .ip(n9266), .ck(clk), .q(
        \pipeline/regfile/data[20][22] ) );
  dp_1 \pipeline/regfile/data_reg[20][23]  ( .ip(n9265), .ck(clk), .q(
        \pipeline/regfile/data[20][23] ) );
  dp_1 \pipeline/regfile/data_reg[20][24]  ( .ip(n9264), .ck(clk), .q(
        \pipeline/regfile/data[20][24] ) );
  dp_1 \pipeline/regfile/data_reg[20][25]  ( .ip(n9263), .ck(clk), .q(
        \pipeline/regfile/data[20][25] ) );
  dp_1 \pipeline/regfile/data_reg[20][26]  ( .ip(n9262), .ck(clk), .q(
        \pipeline/regfile/data[20][26] ) );
  dp_1 \pipeline/regfile/data_reg[20][27]  ( .ip(n9261), .ck(clk), .q(
        \pipeline/regfile/data[20][27] ) );
  dp_1 \pipeline/regfile/data_reg[20][28]  ( .ip(n9260), .ck(clk), .q(
        \pipeline/regfile/data[20][28] ) );
  dp_1 \pipeline/regfile/data_reg[20][29]  ( .ip(n9259), .ck(clk), .q(
        \pipeline/regfile/data[20][29] ) );
  dp_1 \pipeline/regfile/data_reg[20][30]  ( .ip(n9258), .ck(clk), .q(
        \pipeline/regfile/data[20][30] ) );
  dp_1 \pipeline/regfile/data_reg[20][31]  ( .ip(n9257), .ck(clk), .q(
        \pipeline/regfile/data[20][31] ) );
  dp_1 \pipeline/regfile/data_reg[21][0]  ( .ip(n9256), .ck(clk), .q(
        \pipeline/regfile/data[21][0] ) );
  dp_1 \pipeline/regfile/data_reg[21][1]  ( .ip(n9255), .ck(clk), .q(
        \pipeline/regfile/data[21][1] ) );
  dp_1 \pipeline/regfile/data_reg[21][2]  ( .ip(n9254), .ck(clk), .q(
        \pipeline/regfile/data[21][2] ) );
  dp_1 \pipeline/regfile/data_reg[21][3]  ( .ip(n9253), .ck(clk), .q(
        \pipeline/regfile/data[21][3] ) );
  dp_1 \pipeline/regfile/data_reg[21][4]  ( .ip(n9252), .ck(clk), .q(
        \pipeline/regfile/data[21][4] ) );
  dp_1 \pipeline/regfile/data_reg[21][5]  ( .ip(n9251), .ck(clk), .q(
        \pipeline/regfile/data[21][5] ) );
  dp_1 \pipeline/regfile/data_reg[21][6]  ( .ip(n9250), .ck(clk), .q(
        \pipeline/regfile/data[21][6] ) );
  dp_1 \pipeline/regfile/data_reg[21][7]  ( .ip(n9249), .ck(clk), .q(
        \pipeline/regfile/data[21][7] ) );
  dp_1 \pipeline/regfile/data_reg[21][8]  ( .ip(n9248), .ck(clk), .q(
        \pipeline/regfile/data[21][8] ) );
  dp_1 \pipeline/regfile/data_reg[21][9]  ( .ip(n9247), .ck(clk), .q(
        \pipeline/regfile/data[21][9] ) );
  dp_1 \pipeline/regfile/data_reg[21][10]  ( .ip(n9246), .ck(clk), .q(
        \pipeline/regfile/data[21][10] ) );
  dp_1 \pipeline/regfile/data_reg[21][11]  ( .ip(n9245), .ck(clk), .q(
        \pipeline/regfile/data[21][11] ) );
  dp_1 \pipeline/regfile/data_reg[21][12]  ( .ip(n9244), .ck(clk), .q(
        \pipeline/regfile/data[21][12] ) );
  dp_1 \pipeline/regfile/data_reg[21][13]  ( .ip(n9243), .ck(clk), .q(
        \pipeline/regfile/data[21][13] ) );
  dp_1 \pipeline/regfile/data_reg[21][14]  ( .ip(n9242), .ck(clk), .q(
        \pipeline/regfile/data[21][14] ) );
  dp_1 \pipeline/regfile/data_reg[21][15]  ( .ip(n9241), .ck(clk), .q(
        \pipeline/regfile/data[21][15] ) );
  dp_1 \pipeline/regfile/data_reg[21][16]  ( .ip(n9240), .ck(clk), .q(
        \pipeline/regfile/data[21][16] ) );
  dp_1 \pipeline/regfile/data_reg[21][17]  ( .ip(n9239), .ck(clk), .q(
        \pipeline/regfile/data[21][17] ) );
  dp_1 \pipeline/regfile/data_reg[21][18]  ( .ip(n9238), .ck(clk), .q(
        \pipeline/regfile/data[21][18] ) );
  dp_1 \pipeline/regfile/data_reg[21][19]  ( .ip(n9237), .ck(clk), .q(
        \pipeline/regfile/data[21][19] ) );
  dp_1 \pipeline/regfile/data_reg[21][20]  ( .ip(n9236), .ck(clk), .q(
        \pipeline/regfile/data[21][20] ) );
  dp_1 \pipeline/regfile/data_reg[21][21]  ( .ip(n9235), .ck(clk), .q(
        \pipeline/regfile/data[21][21] ) );
  dp_1 \pipeline/regfile/data_reg[21][22]  ( .ip(n9234), .ck(clk), .q(
        \pipeline/regfile/data[21][22] ) );
  dp_1 \pipeline/regfile/data_reg[21][23]  ( .ip(n9233), .ck(clk), .q(
        \pipeline/regfile/data[21][23] ) );
  dp_1 \pipeline/regfile/data_reg[21][24]  ( .ip(n9232), .ck(clk), .q(
        \pipeline/regfile/data[21][24] ) );
  dp_1 \pipeline/regfile/data_reg[21][25]  ( .ip(n9231), .ck(clk), .q(
        \pipeline/regfile/data[21][25] ) );
  dp_1 \pipeline/regfile/data_reg[21][26]  ( .ip(n9230), .ck(clk), .q(
        \pipeline/regfile/data[21][26] ) );
  dp_1 \pipeline/regfile/data_reg[21][27]  ( .ip(n9229), .ck(clk), .q(
        \pipeline/regfile/data[21][27] ) );
  dp_1 \pipeline/regfile/data_reg[21][28]  ( .ip(n9228), .ck(clk), .q(
        \pipeline/regfile/data[21][28] ) );
  dp_1 \pipeline/regfile/data_reg[21][29]  ( .ip(n9227), .ck(clk), .q(
        \pipeline/regfile/data[21][29] ) );
  dp_1 \pipeline/regfile/data_reg[21][30]  ( .ip(n9226), .ck(clk), .q(
        \pipeline/regfile/data[21][30] ) );
  dp_1 \pipeline/regfile/data_reg[21][31]  ( .ip(n9225), .ck(clk), .q(
        \pipeline/regfile/data[21][31] ) );
  dp_1 \pipeline/regfile/data_reg[22][0]  ( .ip(n9224), .ck(clk), .q(
        \pipeline/regfile/data[22][0] ) );
  dp_1 \pipeline/regfile/data_reg[22][1]  ( .ip(n9223), .ck(clk), .q(
        \pipeline/regfile/data[22][1] ) );
  dp_1 \pipeline/regfile/data_reg[22][2]  ( .ip(n9222), .ck(clk), .q(
        \pipeline/regfile/data[22][2] ) );
  dp_1 \pipeline/regfile/data_reg[22][3]  ( .ip(n9221), .ck(clk), .q(
        \pipeline/regfile/data[22][3] ) );
  dp_1 \pipeline/regfile/data_reg[22][4]  ( .ip(n9220), .ck(clk), .q(
        \pipeline/regfile/data[22][4] ) );
  dp_1 \pipeline/regfile/data_reg[22][5]  ( .ip(n9219), .ck(clk), .q(
        \pipeline/regfile/data[22][5] ) );
  dp_1 \pipeline/regfile/data_reg[22][6]  ( .ip(n9218), .ck(clk), .q(
        \pipeline/regfile/data[22][6] ) );
  dp_1 \pipeline/regfile/data_reg[22][7]  ( .ip(n9217), .ck(clk), .q(
        \pipeline/regfile/data[22][7] ) );
  dp_1 \pipeline/regfile/data_reg[22][8]  ( .ip(n9216), .ck(clk), .q(
        \pipeline/regfile/data[22][8] ) );
  dp_1 \pipeline/regfile/data_reg[22][9]  ( .ip(n9215), .ck(clk), .q(
        \pipeline/regfile/data[22][9] ) );
  dp_1 \pipeline/regfile/data_reg[22][10]  ( .ip(n9214), .ck(clk), .q(
        \pipeline/regfile/data[22][10] ) );
  dp_1 \pipeline/regfile/data_reg[22][11]  ( .ip(n9213), .ck(clk), .q(
        \pipeline/regfile/data[22][11] ) );
  dp_1 \pipeline/regfile/data_reg[22][12]  ( .ip(n9212), .ck(clk), .q(
        \pipeline/regfile/data[22][12] ) );
  dp_1 \pipeline/regfile/data_reg[22][13]  ( .ip(n9211), .ck(clk), .q(
        \pipeline/regfile/data[22][13] ) );
  dp_1 \pipeline/regfile/data_reg[22][14]  ( .ip(n9210), .ck(clk), .q(
        \pipeline/regfile/data[22][14] ) );
  dp_1 \pipeline/regfile/data_reg[22][15]  ( .ip(n9209), .ck(clk), .q(
        \pipeline/regfile/data[22][15] ) );
  dp_1 \pipeline/regfile/data_reg[22][16]  ( .ip(n9208), .ck(clk), .q(
        \pipeline/regfile/data[22][16] ) );
  dp_1 \pipeline/regfile/data_reg[22][17]  ( .ip(n9207), .ck(clk), .q(
        \pipeline/regfile/data[22][17] ) );
  dp_1 \pipeline/regfile/data_reg[22][18]  ( .ip(n9206), .ck(clk), .q(
        \pipeline/regfile/data[22][18] ) );
  dp_1 \pipeline/regfile/data_reg[22][19]  ( .ip(n9205), .ck(clk), .q(
        \pipeline/regfile/data[22][19] ) );
  dp_1 \pipeline/regfile/data_reg[22][20]  ( .ip(n9204), .ck(clk), .q(
        \pipeline/regfile/data[22][20] ) );
  dp_1 \pipeline/regfile/data_reg[22][21]  ( .ip(n9203), .ck(clk), .q(
        \pipeline/regfile/data[22][21] ) );
  dp_1 \pipeline/regfile/data_reg[22][22]  ( .ip(n9202), .ck(clk), .q(
        \pipeline/regfile/data[22][22] ) );
  dp_1 \pipeline/regfile/data_reg[22][23]  ( .ip(n9201), .ck(clk), .q(
        \pipeline/regfile/data[22][23] ) );
  dp_1 \pipeline/regfile/data_reg[22][24]  ( .ip(n9200), .ck(clk), .q(
        \pipeline/regfile/data[22][24] ) );
  dp_1 \pipeline/regfile/data_reg[22][25]  ( .ip(n9199), .ck(clk), .q(
        \pipeline/regfile/data[22][25] ) );
  dp_1 \pipeline/regfile/data_reg[22][26]  ( .ip(n9198), .ck(clk), .q(
        \pipeline/regfile/data[22][26] ) );
  dp_1 \pipeline/regfile/data_reg[22][27]  ( .ip(n9197), .ck(clk), .q(
        \pipeline/regfile/data[22][27] ) );
  dp_1 \pipeline/regfile/data_reg[22][28]  ( .ip(n9196), .ck(clk), .q(
        \pipeline/regfile/data[22][28] ) );
  dp_1 \pipeline/regfile/data_reg[22][29]  ( .ip(n9195), .ck(clk), .q(
        \pipeline/regfile/data[22][29] ) );
  dp_1 \pipeline/regfile/data_reg[22][30]  ( .ip(n9194), .ck(clk), .q(
        \pipeline/regfile/data[22][30] ) );
  dp_1 \pipeline/regfile/data_reg[22][31]  ( .ip(n9193), .ck(clk), .q(
        \pipeline/regfile/data[22][31] ) );
  dp_1 \pipeline/regfile/data_reg[23][0]  ( .ip(n9192), .ck(clk), .q(
        \pipeline/regfile/data[23][0] ) );
  dp_1 \pipeline/regfile/data_reg[23][1]  ( .ip(n9191), .ck(clk), .q(
        \pipeline/regfile/data[23][1] ) );
  dp_1 \pipeline/regfile/data_reg[23][2]  ( .ip(n9190), .ck(clk), .q(
        \pipeline/regfile/data[23][2] ) );
  dp_1 \pipeline/regfile/data_reg[23][3]  ( .ip(n9189), .ck(clk), .q(
        \pipeline/regfile/data[23][3] ) );
  dp_1 \pipeline/regfile/data_reg[23][4]  ( .ip(n9188), .ck(clk), .q(
        \pipeline/regfile/data[23][4] ) );
  dp_1 \pipeline/regfile/data_reg[23][5]  ( .ip(n9187), .ck(clk), .q(
        \pipeline/regfile/data[23][5] ) );
  dp_1 \pipeline/regfile/data_reg[23][6]  ( .ip(n9186), .ck(clk), .q(
        \pipeline/regfile/data[23][6] ) );
  dp_1 \pipeline/regfile/data_reg[23][7]  ( .ip(n9185), .ck(clk), .q(
        \pipeline/regfile/data[23][7] ) );
  dp_1 \pipeline/regfile/data_reg[23][8]  ( .ip(n9184), .ck(clk), .q(
        \pipeline/regfile/data[23][8] ) );
  dp_1 \pipeline/regfile/data_reg[23][9]  ( .ip(n9183), .ck(clk), .q(
        \pipeline/regfile/data[23][9] ) );
  dp_1 \pipeline/regfile/data_reg[23][10]  ( .ip(n9182), .ck(clk), .q(
        \pipeline/regfile/data[23][10] ) );
  dp_1 \pipeline/regfile/data_reg[23][11]  ( .ip(n9181), .ck(clk), .q(
        \pipeline/regfile/data[23][11] ) );
  dp_1 \pipeline/regfile/data_reg[23][12]  ( .ip(n9180), .ck(clk), .q(
        \pipeline/regfile/data[23][12] ) );
  dp_1 \pipeline/regfile/data_reg[23][13]  ( .ip(n9179), .ck(clk), .q(
        \pipeline/regfile/data[23][13] ) );
  dp_1 \pipeline/regfile/data_reg[23][14]  ( .ip(n9178), .ck(clk), .q(
        \pipeline/regfile/data[23][14] ) );
  dp_1 \pipeline/regfile/data_reg[23][15]  ( .ip(n9177), .ck(clk), .q(
        \pipeline/regfile/data[23][15] ) );
  dp_1 \pipeline/regfile/data_reg[23][16]  ( .ip(n9176), .ck(clk), .q(
        \pipeline/regfile/data[23][16] ) );
  dp_1 \pipeline/regfile/data_reg[23][17]  ( .ip(n9175), .ck(clk), .q(
        \pipeline/regfile/data[23][17] ) );
  dp_1 \pipeline/regfile/data_reg[23][18]  ( .ip(n9174), .ck(clk), .q(
        \pipeline/regfile/data[23][18] ) );
  dp_1 \pipeline/regfile/data_reg[23][19]  ( .ip(n9173), .ck(clk), .q(
        \pipeline/regfile/data[23][19] ) );
  dp_1 \pipeline/regfile/data_reg[23][20]  ( .ip(n9172), .ck(clk), .q(
        \pipeline/regfile/data[23][20] ) );
  dp_1 \pipeline/regfile/data_reg[23][21]  ( .ip(n9171), .ck(clk), .q(
        \pipeline/regfile/data[23][21] ) );
  dp_1 \pipeline/regfile/data_reg[23][22]  ( .ip(n9170), .ck(clk), .q(
        \pipeline/regfile/data[23][22] ) );
  dp_1 \pipeline/regfile/data_reg[23][23]  ( .ip(n9169), .ck(clk), .q(
        \pipeline/regfile/data[23][23] ) );
  dp_1 \pipeline/regfile/data_reg[23][24]  ( .ip(n9168), .ck(clk), .q(
        \pipeline/regfile/data[23][24] ) );
  dp_1 \pipeline/regfile/data_reg[23][25]  ( .ip(n9167), .ck(clk), .q(
        \pipeline/regfile/data[23][25] ) );
  dp_1 \pipeline/regfile/data_reg[23][26]  ( .ip(n9166), .ck(clk), .q(
        \pipeline/regfile/data[23][26] ) );
  dp_1 \pipeline/regfile/data_reg[23][27]  ( .ip(n9165), .ck(clk), .q(
        \pipeline/regfile/data[23][27] ) );
  dp_1 \pipeline/regfile/data_reg[23][28]  ( .ip(n9164), .ck(clk), .q(
        \pipeline/regfile/data[23][28] ) );
  dp_1 \pipeline/regfile/data_reg[23][29]  ( .ip(n9163), .ck(clk), .q(
        \pipeline/regfile/data[23][29] ) );
  dp_1 \pipeline/regfile/data_reg[23][30]  ( .ip(n9162), .ck(clk), .q(
        \pipeline/regfile/data[23][30] ) );
  dp_1 \pipeline/regfile/data_reg[23][31]  ( .ip(n9161), .ck(clk), .q(
        \pipeline/regfile/data[23][31] ) );
  dp_1 \pipeline/regfile/data_reg[24][0]  ( .ip(n9160), .ck(clk), .q(
        \pipeline/regfile/data[24][0] ) );
  dp_1 \pipeline/regfile/data_reg[24][1]  ( .ip(n9159), .ck(clk), .q(
        \pipeline/regfile/data[24][1] ) );
  dp_1 \pipeline/regfile/data_reg[24][2]  ( .ip(n9158), .ck(clk), .q(
        \pipeline/regfile/data[24][2] ) );
  dp_1 \pipeline/regfile/data_reg[24][3]  ( .ip(n9157), .ck(clk), .q(
        \pipeline/regfile/data[24][3] ) );
  dp_1 \pipeline/regfile/data_reg[24][4]  ( .ip(n9156), .ck(clk), .q(
        \pipeline/regfile/data[24][4] ) );
  dp_1 \pipeline/regfile/data_reg[24][5]  ( .ip(n9155), .ck(clk), .q(
        \pipeline/regfile/data[24][5] ) );
  dp_1 \pipeline/regfile/data_reg[24][6]  ( .ip(n9154), .ck(clk), .q(
        \pipeline/regfile/data[24][6] ) );
  dp_1 \pipeline/regfile/data_reg[24][7]  ( .ip(n9153), .ck(clk), .q(
        \pipeline/regfile/data[24][7] ) );
  dp_1 \pipeline/regfile/data_reg[24][8]  ( .ip(n9152), .ck(clk), .q(
        \pipeline/regfile/data[24][8] ) );
  dp_1 \pipeline/regfile/data_reg[24][9]  ( .ip(n9151), .ck(clk), .q(
        \pipeline/regfile/data[24][9] ) );
  dp_1 \pipeline/regfile/data_reg[24][10]  ( .ip(n9150), .ck(clk), .q(
        \pipeline/regfile/data[24][10] ) );
  dp_1 \pipeline/regfile/data_reg[24][11]  ( .ip(n9149), .ck(clk), .q(
        \pipeline/regfile/data[24][11] ) );
  dp_1 \pipeline/regfile/data_reg[24][12]  ( .ip(n9148), .ck(clk), .q(
        \pipeline/regfile/data[24][12] ) );
  dp_1 \pipeline/regfile/data_reg[24][13]  ( .ip(n9147), .ck(clk), .q(
        \pipeline/regfile/data[24][13] ) );
  dp_1 \pipeline/regfile/data_reg[24][14]  ( .ip(n9146), .ck(clk), .q(
        \pipeline/regfile/data[24][14] ) );
  dp_1 \pipeline/regfile/data_reg[24][15]  ( .ip(n9145), .ck(clk), .q(
        \pipeline/regfile/data[24][15] ) );
  dp_1 \pipeline/regfile/data_reg[24][16]  ( .ip(n9144), .ck(clk), .q(
        \pipeline/regfile/data[24][16] ) );
  dp_1 \pipeline/regfile/data_reg[24][17]  ( .ip(n9143), .ck(clk), .q(
        \pipeline/regfile/data[24][17] ) );
  dp_1 \pipeline/regfile/data_reg[24][18]  ( .ip(n9142), .ck(clk), .q(
        \pipeline/regfile/data[24][18] ) );
  dp_1 \pipeline/regfile/data_reg[24][19]  ( .ip(n9141), .ck(clk), .q(
        \pipeline/regfile/data[24][19] ) );
  dp_1 \pipeline/regfile/data_reg[24][20]  ( .ip(n9140), .ck(clk), .q(
        \pipeline/regfile/data[24][20] ) );
  dp_1 \pipeline/regfile/data_reg[24][21]  ( .ip(n9139), .ck(clk), .q(
        \pipeline/regfile/data[24][21] ) );
  dp_1 \pipeline/regfile/data_reg[24][22]  ( .ip(n9138), .ck(clk), .q(
        \pipeline/regfile/data[24][22] ) );
  dp_1 \pipeline/regfile/data_reg[24][23]  ( .ip(n9137), .ck(clk), .q(
        \pipeline/regfile/data[24][23] ) );
  dp_1 \pipeline/regfile/data_reg[24][24]  ( .ip(n9136), .ck(clk), .q(
        \pipeline/regfile/data[24][24] ) );
  dp_1 \pipeline/regfile/data_reg[24][25]  ( .ip(n9135), .ck(clk), .q(
        \pipeline/regfile/data[24][25] ) );
  dp_1 \pipeline/regfile/data_reg[24][26]  ( .ip(n9134), .ck(clk), .q(
        \pipeline/regfile/data[24][26] ) );
  dp_1 \pipeline/regfile/data_reg[24][27]  ( .ip(n9133), .ck(clk), .q(
        \pipeline/regfile/data[24][27] ) );
  dp_1 \pipeline/regfile/data_reg[24][28]  ( .ip(n9132), .ck(clk), .q(
        \pipeline/regfile/data[24][28] ) );
  dp_1 \pipeline/regfile/data_reg[24][29]  ( .ip(n9131), .ck(clk), .q(
        \pipeline/regfile/data[24][29] ) );
  dp_1 \pipeline/regfile/data_reg[24][30]  ( .ip(n9130), .ck(clk), .q(
        \pipeline/regfile/data[24][30] ) );
  dp_1 \pipeline/regfile/data_reg[24][31]  ( .ip(n9129), .ck(clk), .q(
        \pipeline/regfile/data[24][31] ) );
  dp_1 \pipeline/regfile/data_reg[25][0]  ( .ip(n9128), .ck(clk), .q(
        \pipeline/regfile/data[25][0] ) );
  dp_1 \pipeline/regfile/data_reg[25][1]  ( .ip(n9127), .ck(clk), .q(
        \pipeline/regfile/data[25][1] ) );
  dp_1 \pipeline/regfile/data_reg[25][2]  ( .ip(n9126), .ck(clk), .q(
        \pipeline/regfile/data[25][2] ) );
  dp_1 \pipeline/regfile/data_reg[25][3]  ( .ip(n9125), .ck(clk), .q(
        \pipeline/regfile/data[25][3] ) );
  dp_1 \pipeline/regfile/data_reg[25][4]  ( .ip(n9124), .ck(clk), .q(
        \pipeline/regfile/data[25][4] ) );
  dp_1 \pipeline/regfile/data_reg[25][5]  ( .ip(n9123), .ck(clk), .q(
        \pipeline/regfile/data[25][5] ) );
  dp_1 \pipeline/regfile/data_reg[25][6]  ( .ip(n9122), .ck(clk), .q(
        \pipeline/regfile/data[25][6] ) );
  dp_1 \pipeline/regfile/data_reg[25][7]  ( .ip(n9121), .ck(clk), .q(
        \pipeline/regfile/data[25][7] ) );
  dp_1 \pipeline/regfile/data_reg[25][8]  ( .ip(n9120), .ck(clk), .q(
        \pipeline/regfile/data[25][8] ) );
  dp_1 \pipeline/regfile/data_reg[25][9]  ( .ip(n9119), .ck(clk), .q(
        \pipeline/regfile/data[25][9] ) );
  dp_1 \pipeline/regfile/data_reg[25][10]  ( .ip(n9118), .ck(clk), .q(
        \pipeline/regfile/data[25][10] ) );
  dp_1 \pipeline/regfile/data_reg[25][11]  ( .ip(n9117), .ck(clk), .q(
        \pipeline/regfile/data[25][11] ) );
  dp_1 \pipeline/regfile/data_reg[25][12]  ( .ip(n9116), .ck(clk), .q(
        \pipeline/regfile/data[25][12] ) );
  dp_1 \pipeline/regfile/data_reg[25][13]  ( .ip(n9115), .ck(clk), .q(
        \pipeline/regfile/data[25][13] ) );
  dp_1 \pipeline/regfile/data_reg[25][14]  ( .ip(n9114), .ck(clk), .q(
        \pipeline/regfile/data[25][14] ) );
  dp_1 \pipeline/regfile/data_reg[25][15]  ( .ip(n9113), .ck(clk), .q(
        \pipeline/regfile/data[25][15] ) );
  dp_1 \pipeline/regfile/data_reg[25][16]  ( .ip(n9112), .ck(clk), .q(
        \pipeline/regfile/data[25][16] ) );
  dp_1 \pipeline/regfile/data_reg[25][17]  ( .ip(n9111), .ck(clk), .q(
        \pipeline/regfile/data[25][17] ) );
  dp_1 \pipeline/regfile/data_reg[25][18]  ( .ip(n9110), .ck(clk), .q(
        \pipeline/regfile/data[25][18] ) );
  dp_1 \pipeline/regfile/data_reg[25][19]  ( .ip(n9109), .ck(clk), .q(
        \pipeline/regfile/data[25][19] ) );
  dp_1 \pipeline/regfile/data_reg[25][20]  ( .ip(n9108), .ck(clk), .q(
        \pipeline/regfile/data[25][20] ) );
  dp_1 \pipeline/regfile/data_reg[25][21]  ( .ip(n9107), .ck(clk), .q(
        \pipeline/regfile/data[25][21] ) );
  dp_1 \pipeline/regfile/data_reg[25][22]  ( .ip(n9106), .ck(clk), .q(
        \pipeline/regfile/data[25][22] ) );
  dp_1 \pipeline/regfile/data_reg[25][23]  ( .ip(n9105), .ck(clk), .q(
        \pipeline/regfile/data[25][23] ) );
  dp_1 \pipeline/regfile/data_reg[25][24]  ( .ip(n9104), .ck(clk), .q(
        \pipeline/regfile/data[25][24] ) );
  dp_1 \pipeline/regfile/data_reg[25][25]  ( .ip(n9103), .ck(clk), .q(
        \pipeline/regfile/data[25][25] ) );
  dp_1 \pipeline/regfile/data_reg[25][26]  ( .ip(n9102), .ck(clk), .q(
        \pipeline/regfile/data[25][26] ) );
  dp_1 \pipeline/regfile/data_reg[25][27]  ( .ip(n9101), .ck(clk), .q(
        \pipeline/regfile/data[25][27] ) );
  dp_1 \pipeline/regfile/data_reg[25][28]  ( .ip(n9100), .ck(clk), .q(
        \pipeline/regfile/data[25][28] ) );
  dp_1 \pipeline/regfile/data_reg[25][29]  ( .ip(n9099), .ck(clk), .q(
        \pipeline/regfile/data[25][29] ) );
  dp_1 \pipeline/regfile/data_reg[25][30]  ( .ip(n9098), .ck(clk), .q(
        \pipeline/regfile/data[25][30] ) );
  dp_1 \pipeline/regfile/data_reg[25][31]  ( .ip(n9097), .ck(clk), .q(
        \pipeline/regfile/data[25][31] ) );
  dp_1 \pipeline/regfile/data_reg[26][0]  ( .ip(n9096), .ck(clk), .q(
        \pipeline/regfile/data[26][0] ) );
  dp_1 \pipeline/regfile/data_reg[26][1]  ( .ip(n9095), .ck(clk), .q(
        \pipeline/regfile/data[26][1] ) );
  dp_1 \pipeline/regfile/data_reg[26][2]  ( .ip(n9094), .ck(clk), .q(
        \pipeline/regfile/data[26][2] ) );
  dp_1 \pipeline/regfile/data_reg[26][3]  ( .ip(n9093), .ck(clk), .q(
        \pipeline/regfile/data[26][3] ) );
  dp_1 \pipeline/regfile/data_reg[26][4]  ( .ip(n9092), .ck(clk), .q(
        \pipeline/regfile/data[26][4] ) );
  dp_1 \pipeline/regfile/data_reg[26][5]  ( .ip(n9091), .ck(clk), .q(
        \pipeline/regfile/data[26][5] ) );
  dp_1 \pipeline/regfile/data_reg[26][6]  ( .ip(n9090), .ck(clk), .q(
        \pipeline/regfile/data[26][6] ) );
  dp_1 \pipeline/regfile/data_reg[26][7]  ( .ip(n9089), .ck(clk), .q(
        \pipeline/regfile/data[26][7] ) );
  dp_1 \pipeline/regfile/data_reg[26][8]  ( .ip(n9088), .ck(clk), .q(
        \pipeline/regfile/data[26][8] ) );
  dp_1 \pipeline/regfile/data_reg[26][9]  ( .ip(n9087), .ck(clk), .q(
        \pipeline/regfile/data[26][9] ) );
  dp_1 \pipeline/regfile/data_reg[26][10]  ( .ip(n9086), .ck(clk), .q(
        \pipeline/regfile/data[26][10] ) );
  dp_1 \pipeline/regfile/data_reg[26][11]  ( .ip(n9085), .ck(clk), .q(
        \pipeline/regfile/data[26][11] ) );
  dp_1 \pipeline/regfile/data_reg[26][12]  ( .ip(n9084), .ck(clk), .q(
        \pipeline/regfile/data[26][12] ) );
  dp_1 \pipeline/regfile/data_reg[26][13]  ( .ip(n9083), .ck(clk), .q(
        \pipeline/regfile/data[26][13] ) );
  dp_1 \pipeline/regfile/data_reg[26][14]  ( .ip(n9082), .ck(clk), .q(
        \pipeline/regfile/data[26][14] ) );
  dp_1 \pipeline/regfile/data_reg[26][15]  ( .ip(n9081), .ck(clk), .q(
        \pipeline/regfile/data[26][15] ) );
  dp_1 \pipeline/regfile/data_reg[26][16]  ( .ip(n9080), .ck(clk), .q(
        \pipeline/regfile/data[26][16] ) );
  dp_1 \pipeline/regfile/data_reg[26][17]  ( .ip(n9079), .ck(clk), .q(
        \pipeline/regfile/data[26][17] ) );
  dp_1 \pipeline/regfile/data_reg[26][18]  ( .ip(n9078), .ck(clk), .q(
        \pipeline/regfile/data[26][18] ) );
  dp_1 \pipeline/regfile/data_reg[26][19]  ( .ip(n9077), .ck(clk), .q(
        \pipeline/regfile/data[26][19] ) );
  dp_1 \pipeline/regfile/data_reg[26][20]  ( .ip(n9076), .ck(clk), .q(
        \pipeline/regfile/data[26][20] ) );
  dp_1 \pipeline/regfile/data_reg[26][21]  ( .ip(n9075), .ck(clk), .q(
        \pipeline/regfile/data[26][21] ) );
  dp_1 \pipeline/regfile/data_reg[26][22]  ( .ip(n9074), .ck(clk), .q(
        \pipeline/regfile/data[26][22] ) );
  dp_1 \pipeline/regfile/data_reg[26][23]  ( .ip(n9073), .ck(clk), .q(
        \pipeline/regfile/data[26][23] ) );
  dp_1 \pipeline/regfile/data_reg[26][24]  ( .ip(n9072), .ck(clk), .q(
        \pipeline/regfile/data[26][24] ) );
  dp_1 \pipeline/regfile/data_reg[26][25]  ( .ip(n9071), .ck(clk), .q(
        \pipeline/regfile/data[26][25] ) );
  dp_1 \pipeline/regfile/data_reg[26][26]  ( .ip(n9070), .ck(clk), .q(
        \pipeline/regfile/data[26][26] ) );
  dp_1 \pipeline/regfile/data_reg[26][27]  ( .ip(n9069), .ck(clk), .q(
        \pipeline/regfile/data[26][27] ) );
  dp_1 \pipeline/regfile/data_reg[26][28]  ( .ip(n9068), .ck(clk), .q(
        \pipeline/regfile/data[26][28] ) );
  dp_1 \pipeline/regfile/data_reg[26][29]  ( .ip(n9067), .ck(clk), .q(
        \pipeline/regfile/data[26][29] ) );
  dp_1 \pipeline/regfile/data_reg[26][30]  ( .ip(n9066), .ck(clk), .q(
        \pipeline/regfile/data[26][30] ) );
  dp_1 \pipeline/regfile/data_reg[26][31]  ( .ip(n9065), .ck(clk), .q(
        \pipeline/regfile/data[26][31] ) );
  dp_1 \pipeline/regfile/data_reg[27][0]  ( .ip(n9064), .ck(clk), .q(
        \pipeline/regfile/data[27][0] ) );
  dp_1 \pipeline/regfile/data_reg[27][1]  ( .ip(n9063), .ck(clk), .q(
        \pipeline/regfile/data[27][1] ) );
  dp_1 \pipeline/regfile/data_reg[27][2]  ( .ip(n9062), .ck(clk), .q(
        \pipeline/regfile/data[27][2] ) );
  dp_1 \pipeline/regfile/data_reg[27][3]  ( .ip(n9061), .ck(clk), .q(
        \pipeline/regfile/data[27][3] ) );
  dp_1 \pipeline/regfile/data_reg[27][4]  ( .ip(n9060), .ck(clk), .q(
        \pipeline/regfile/data[27][4] ) );
  dp_1 \pipeline/regfile/data_reg[27][5]  ( .ip(n9059), .ck(clk), .q(
        \pipeline/regfile/data[27][5] ) );
  dp_1 \pipeline/regfile/data_reg[27][6]  ( .ip(n9058), .ck(clk), .q(
        \pipeline/regfile/data[27][6] ) );
  dp_1 \pipeline/regfile/data_reg[27][7]  ( .ip(n9057), .ck(clk), .q(
        \pipeline/regfile/data[27][7] ) );
  dp_1 \pipeline/regfile/data_reg[27][8]  ( .ip(n9056), .ck(clk), .q(
        \pipeline/regfile/data[27][8] ) );
  dp_1 \pipeline/regfile/data_reg[27][9]  ( .ip(n9055), .ck(clk), .q(
        \pipeline/regfile/data[27][9] ) );
  dp_1 \pipeline/regfile/data_reg[27][10]  ( .ip(n9054), .ck(clk), .q(
        \pipeline/regfile/data[27][10] ) );
  dp_1 \pipeline/regfile/data_reg[27][11]  ( .ip(n9053), .ck(clk), .q(
        \pipeline/regfile/data[27][11] ) );
  dp_1 \pipeline/regfile/data_reg[27][12]  ( .ip(n9052), .ck(clk), .q(
        \pipeline/regfile/data[27][12] ) );
  dp_1 \pipeline/regfile/data_reg[27][13]  ( .ip(n9051), .ck(clk), .q(
        \pipeline/regfile/data[27][13] ) );
  dp_1 \pipeline/regfile/data_reg[27][14]  ( .ip(n9050), .ck(clk), .q(
        \pipeline/regfile/data[27][14] ) );
  dp_1 \pipeline/regfile/data_reg[27][15]  ( .ip(n9049), .ck(clk), .q(
        \pipeline/regfile/data[27][15] ) );
  dp_1 \pipeline/regfile/data_reg[27][16]  ( .ip(n9048), .ck(clk), .q(
        \pipeline/regfile/data[27][16] ) );
  dp_1 \pipeline/regfile/data_reg[27][17]  ( .ip(n9047), .ck(clk), .q(
        \pipeline/regfile/data[27][17] ) );
  dp_1 \pipeline/regfile/data_reg[27][18]  ( .ip(n9046), .ck(clk), .q(
        \pipeline/regfile/data[27][18] ) );
  dp_1 \pipeline/regfile/data_reg[27][19]  ( .ip(n9045), .ck(clk), .q(
        \pipeline/regfile/data[27][19] ) );
  dp_1 \pipeline/regfile/data_reg[27][20]  ( .ip(n9044), .ck(clk), .q(
        \pipeline/regfile/data[27][20] ) );
  dp_1 \pipeline/regfile/data_reg[27][21]  ( .ip(n9043), .ck(clk), .q(
        \pipeline/regfile/data[27][21] ) );
  dp_1 \pipeline/regfile/data_reg[27][22]  ( .ip(n9042), .ck(clk), .q(
        \pipeline/regfile/data[27][22] ) );
  dp_1 \pipeline/regfile/data_reg[27][23]  ( .ip(n9041), .ck(clk), .q(
        \pipeline/regfile/data[27][23] ) );
  dp_1 \pipeline/regfile/data_reg[27][24]  ( .ip(n9040), .ck(clk), .q(
        \pipeline/regfile/data[27][24] ) );
  dp_1 \pipeline/regfile/data_reg[27][25]  ( .ip(n9039), .ck(clk), .q(
        \pipeline/regfile/data[27][25] ) );
  dp_1 \pipeline/regfile/data_reg[27][26]  ( .ip(n9038), .ck(clk), .q(
        \pipeline/regfile/data[27][26] ) );
  dp_1 \pipeline/regfile/data_reg[27][27]  ( .ip(n9037), .ck(clk), .q(
        \pipeline/regfile/data[27][27] ) );
  dp_1 \pipeline/regfile/data_reg[27][28]  ( .ip(n9036), .ck(clk), .q(
        \pipeline/regfile/data[27][28] ) );
  dp_1 \pipeline/regfile/data_reg[27][29]  ( .ip(n9035), .ck(clk), .q(
        \pipeline/regfile/data[27][29] ) );
  dp_1 \pipeline/regfile/data_reg[27][30]  ( .ip(n9034), .ck(clk), .q(
        \pipeline/regfile/data[27][30] ) );
  dp_1 \pipeline/regfile/data_reg[27][31]  ( .ip(n9033), .ck(clk), .q(
        \pipeline/regfile/data[27][31] ) );
  dp_1 \pipeline/regfile/data_reg[28][0]  ( .ip(n9032), .ck(clk), .q(
        \pipeline/regfile/data[28][0] ) );
  dp_1 \pipeline/regfile/data_reg[28][1]  ( .ip(n9031), .ck(clk), .q(
        \pipeline/regfile/data[28][1] ) );
  dp_1 \pipeline/regfile/data_reg[28][2]  ( .ip(n9030), .ck(clk), .q(
        \pipeline/regfile/data[28][2] ) );
  dp_1 \pipeline/regfile/data_reg[28][3]  ( .ip(n9029), .ck(clk), .q(
        \pipeline/regfile/data[28][3] ) );
  dp_1 \pipeline/regfile/data_reg[28][4]  ( .ip(n9028), .ck(clk), .q(
        \pipeline/regfile/data[28][4] ) );
  dp_1 \pipeline/regfile/data_reg[28][5]  ( .ip(n9027), .ck(clk), .q(
        \pipeline/regfile/data[28][5] ) );
  dp_1 \pipeline/regfile/data_reg[28][6]  ( .ip(n9026), .ck(clk), .q(
        \pipeline/regfile/data[28][6] ) );
  dp_1 \pipeline/regfile/data_reg[28][7]  ( .ip(n9025), .ck(clk), .q(
        \pipeline/regfile/data[28][7] ) );
  dp_1 \pipeline/regfile/data_reg[28][8]  ( .ip(n9024), .ck(clk), .q(
        \pipeline/regfile/data[28][8] ) );
  dp_1 \pipeline/regfile/data_reg[28][9]  ( .ip(n9023), .ck(clk), .q(
        \pipeline/regfile/data[28][9] ) );
  dp_1 \pipeline/regfile/data_reg[28][10]  ( .ip(n9022), .ck(clk), .q(
        \pipeline/regfile/data[28][10] ) );
  dp_1 \pipeline/regfile/data_reg[28][11]  ( .ip(n9021), .ck(clk), .q(
        \pipeline/regfile/data[28][11] ) );
  dp_1 \pipeline/regfile/data_reg[28][12]  ( .ip(n9020), .ck(clk), .q(
        \pipeline/regfile/data[28][12] ) );
  dp_1 \pipeline/regfile/data_reg[28][13]  ( .ip(n9019), .ck(clk), .q(
        \pipeline/regfile/data[28][13] ) );
  dp_1 \pipeline/regfile/data_reg[28][14]  ( .ip(n9018), .ck(clk), .q(
        \pipeline/regfile/data[28][14] ) );
  dp_1 \pipeline/regfile/data_reg[28][15]  ( .ip(n9017), .ck(clk), .q(
        \pipeline/regfile/data[28][15] ) );
  dp_1 \pipeline/regfile/data_reg[28][16]  ( .ip(n9016), .ck(clk), .q(
        \pipeline/regfile/data[28][16] ) );
  dp_1 \pipeline/regfile/data_reg[28][17]  ( .ip(n9015), .ck(clk), .q(
        \pipeline/regfile/data[28][17] ) );
  dp_1 \pipeline/regfile/data_reg[28][18]  ( .ip(n9014), .ck(clk), .q(
        \pipeline/regfile/data[28][18] ) );
  dp_1 \pipeline/regfile/data_reg[28][19]  ( .ip(n9013), .ck(clk), .q(
        \pipeline/regfile/data[28][19] ) );
  dp_1 \pipeline/regfile/data_reg[28][20]  ( .ip(n9012), .ck(clk), .q(
        \pipeline/regfile/data[28][20] ) );
  dp_1 \pipeline/regfile/data_reg[28][21]  ( .ip(n9011), .ck(clk), .q(
        \pipeline/regfile/data[28][21] ) );
  dp_1 \pipeline/regfile/data_reg[28][22]  ( .ip(n9010), .ck(clk), .q(
        \pipeline/regfile/data[28][22] ) );
  dp_1 \pipeline/regfile/data_reg[28][23]  ( .ip(n9009), .ck(clk), .q(
        \pipeline/regfile/data[28][23] ) );
  dp_1 \pipeline/regfile/data_reg[28][24]  ( .ip(n9008), .ck(clk), .q(
        \pipeline/regfile/data[28][24] ) );
  dp_1 \pipeline/regfile/data_reg[28][25]  ( .ip(n9007), .ck(clk), .q(
        \pipeline/regfile/data[28][25] ) );
  dp_1 \pipeline/regfile/data_reg[28][26]  ( .ip(n9006), .ck(clk), .q(
        \pipeline/regfile/data[28][26] ) );
  dp_1 \pipeline/regfile/data_reg[28][27]  ( .ip(n9005), .ck(clk), .q(
        \pipeline/regfile/data[28][27] ) );
  dp_1 \pipeline/regfile/data_reg[28][28]  ( .ip(n9004), .ck(clk), .q(
        \pipeline/regfile/data[28][28] ) );
  dp_1 \pipeline/regfile/data_reg[28][29]  ( .ip(n9003), .ck(clk), .q(
        \pipeline/regfile/data[28][29] ) );
  dp_1 \pipeline/regfile/data_reg[28][30]  ( .ip(n9002), .ck(clk), .q(
        \pipeline/regfile/data[28][30] ) );
  dp_1 \pipeline/regfile/data_reg[28][31]  ( .ip(n9001), .ck(clk), .q(
        \pipeline/regfile/data[28][31] ) );
  dp_1 \pipeline/regfile/data_reg[29][0]  ( .ip(n9000), .ck(clk), .q(
        \pipeline/regfile/data[29][0] ) );
  dp_1 \pipeline/regfile/data_reg[29][1]  ( .ip(n8999), .ck(clk), .q(
        \pipeline/regfile/data[29][1] ) );
  dp_1 \pipeline/regfile/data_reg[29][2]  ( .ip(n8998), .ck(clk), .q(
        \pipeline/regfile/data[29][2] ) );
  dp_1 \pipeline/regfile/data_reg[29][3]  ( .ip(n8997), .ck(clk), .q(
        \pipeline/regfile/data[29][3] ) );
  dp_1 \pipeline/regfile/data_reg[29][4]  ( .ip(n8996), .ck(clk), .q(
        \pipeline/regfile/data[29][4] ) );
  dp_1 \pipeline/regfile/data_reg[29][5]  ( .ip(n8995), .ck(clk), .q(
        \pipeline/regfile/data[29][5] ) );
  dp_1 \pipeline/regfile/data_reg[29][6]  ( .ip(n8994), .ck(clk), .q(
        \pipeline/regfile/data[29][6] ) );
  dp_1 \pipeline/regfile/data_reg[29][7]  ( .ip(n8993), .ck(clk), .q(
        \pipeline/regfile/data[29][7] ) );
  dp_1 \pipeline/regfile/data_reg[29][8]  ( .ip(n8992), .ck(clk), .q(
        \pipeline/regfile/data[29][8] ) );
  dp_1 \pipeline/regfile/data_reg[29][9]  ( .ip(n8991), .ck(clk), .q(
        \pipeline/regfile/data[29][9] ) );
  dp_1 \pipeline/regfile/data_reg[29][10]  ( .ip(n8990), .ck(clk), .q(
        \pipeline/regfile/data[29][10] ) );
  dp_1 \pipeline/regfile/data_reg[29][11]  ( .ip(n8989), .ck(clk), .q(
        \pipeline/regfile/data[29][11] ) );
  dp_1 \pipeline/regfile/data_reg[29][12]  ( .ip(n8988), .ck(clk), .q(
        \pipeline/regfile/data[29][12] ) );
  dp_1 \pipeline/regfile/data_reg[29][13]  ( .ip(n8987), .ck(clk), .q(
        \pipeline/regfile/data[29][13] ) );
  dp_1 \pipeline/regfile/data_reg[29][14]  ( .ip(n8986), .ck(clk), .q(
        \pipeline/regfile/data[29][14] ) );
  dp_1 \pipeline/regfile/data_reg[29][15]  ( .ip(n8985), .ck(clk), .q(
        \pipeline/regfile/data[29][15] ) );
  dp_1 \pipeline/regfile/data_reg[29][16]  ( .ip(n8984), .ck(clk), .q(
        \pipeline/regfile/data[29][16] ) );
  dp_1 \pipeline/regfile/data_reg[29][17]  ( .ip(n8983), .ck(clk), .q(
        \pipeline/regfile/data[29][17] ) );
  dp_1 \pipeline/regfile/data_reg[29][18]  ( .ip(n8982), .ck(clk), .q(
        \pipeline/regfile/data[29][18] ) );
  dp_1 \pipeline/regfile/data_reg[29][19]  ( .ip(n8981), .ck(clk), .q(
        \pipeline/regfile/data[29][19] ) );
  dp_1 \pipeline/regfile/data_reg[29][20]  ( .ip(n8980), .ck(clk), .q(
        \pipeline/regfile/data[29][20] ) );
  dp_1 \pipeline/regfile/data_reg[29][21]  ( .ip(n8979), .ck(clk), .q(
        \pipeline/regfile/data[29][21] ) );
  dp_1 \pipeline/regfile/data_reg[29][22]  ( .ip(n8978), .ck(clk), .q(
        \pipeline/regfile/data[29][22] ) );
  dp_1 \pipeline/regfile/data_reg[29][23]  ( .ip(n8977), .ck(clk), .q(
        \pipeline/regfile/data[29][23] ) );
  dp_1 \pipeline/regfile/data_reg[29][24]  ( .ip(n8976), .ck(clk), .q(
        \pipeline/regfile/data[29][24] ) );
  dp_1 \pipeline/regfile/data_reg[29][25]  ( .ip(n8975), .ck(clk), .q(
        \pipeline/regfile/data[29][25] ) );
  dp_1 \pipeline/regfile/data_reg[29][26]  ( .ip(n8974), .ck(clk), .q(
        \pipeline/regfile/data[29][26] ) );
  dp_1 \pipeline/regfile/data_reg[29][27]  ( .ip(n8973), .ck(clk), .q(
        \pipeline/regfile/data[29][27] ) );
  dp_1 \pipeline/regfile/data_reg[29][28]  ( .ip(n8972), .ck(clk), .q(
        \pipeline/regfile/data[29][28] ) );
  dp_1 \pipeline/regfile/data_reg[29][29]  ( .ip(n8971), .ck(clk), .q(
        \pipeline/regfile/data[29][29] ) );
  dp_1 \pipeline/regfile/data_reg[29][30]  ( .ip(n8970), .ck(clk), .q(
        \pipeline/regfile/data[29][30] ) );
  dp_1 \pipeline/regfile/data_reg[29][31]  ( .ip(n8969), .ck(clk), .q(
        \pipeline/regfile/data[29][31] ) );
  dp_1 \pipeline/regfile/data_reg[30][0]  ( .ip(n8968), .ck(clk), .q(
        \pipeline/regfile/data[30][0] ) );
  dp_1 \pipeline/regfile/data_reg[30][1]  ( .ip(n8967), .ck(clk), .q(
        \pipeline/regfile/data[30][1] ) );
  dp_1 \pipeline/regfile/data_reg[30][2]  ( .ip(n8966), .ck(clk), .q(
        \pipeline/regfile/data[30][2] ) );
  dp_1 \pipeline/regfile/data_reg[30][3]  ( .ip(n8965), .ck(clk), .q(
        \pipeline/regfile/data[30][3] ) );
  dp_1 \pipeline/regfile/data_reg[30][4]  ( .ip(n8964), .ck(clk), .q(
        \pipeline/regfile/data[30][4] ) );
  dp_1 \pipeline/regfile/data_reg[30][5]  ( .ip(n8963), .ck(clk), .q(
        \pipeline/regfile/data[30][5] ) );
  dp_1 \pipeline/regfile/data_reg[30][6]  ( .ip(n8962), .ck(clk), .q(
        \pipeline/regfile/data[30][6] ) );
  dp_1 \pipeline/regfile/data_reg[30][7]  ( .ip(n8961), .ck(clk), .q(
        \pipeline/regfile/data[30][7] ) );
  dp_1 \pipeline/regfile/data_reg[30][8]  ( .ip(n8960), .ck(clk), .q(
        \pipeline/regfile/data[30][8] ) );
  dp_1 \pipeline/regfile/data_reg[30][9]  ( .ip(n8959), .ck(clk), .q(
        \pipeline/regfile/data[30][9] ) );
  dp_1 \pipeline/regfile/data_reg[30][10]  ( .ip(n8958), .ck(clk), .q(
        \pipeline/regfile/data[30][10] ) );
  dp_1 \pipeline/regfile/data_reg[30][11]  ( .ip(n8957), .ck(clk), .q(
        \pipeline/regfile/data[30][11] ) );
  dp_1 \pipeline/regfile/data_reg[30][12]  ( .ip(n8956), .ck(clk), .q(
        \pipeline/regfile/data[30][12] ) );
  dp_1 \pipeline/regfile/data_reg[30][13]  ( .ip(n8955), .ck(clk), .q(
        \pipeline/regfile/data[30][13] ) );
  dp_1 \pipeline/regfile/data_reg[30][14]  ( .ip(n8954), .ck(clk), .q(
        \pipeline/regfile/data[30][14] ) );
  dp_1 \pipeline/regfile/data_reg[30][15]  ( .ip(n8953), .ck(clk), .q(
        \pipeline/regfile/data[30][15] ) );
  dp_1 \pipeline/regfile/data_reg[30][16]  ( .ip(n8952), .ck(clk), .q(
        \pipeline/regfile/data[30][16] ) );
  dp_1 \pipeline/regfile/data_reg[30][17]  ( .ip(n8951), .ck(clk), .q(
        \pipeline/regfile/data[30][17] ) );
  dp_1 \pipeline/regfile/data_reg[30][18]  ( .ip(n8950), .ck(clk), .q(
        \pipeline/regfile/data[30][18] ) );
  dp_1 \pipeline/regfile/data_reg[30][19]  ( .ip(n8949), .ck(clk), .q(
        \pipeline/regfile/data[30][19] ) );
  dp_1 \pipeline/regfile/data_reg[30][20]  ( .ip(n8948), .ck(clk), .q(
        \pipeline/regfile/data[30][20] ) );
  dp_1 \pipeline/regfile/data_reg[30][21]  ( .ip(n8947), .ck(clk), .q(
        \pipeline/regfile/data[30][21] ) );
  dp_1 \pipeline/regfile/data_reg[30][22]  ( .ip(n8946), .ck(clk), .q(
        \pipeline/regfile/data[30][22] ) );
  dp_1 \pipeline/regfile/data_reg[30][23]  ( .ip(n8945), .ck(clk), .q(
        \pipeline/regfile/data[30][23] ) );
  dp_1 \pipeline/regfile/data_reg[30][24]  ( .ip(n8944), .ck(clk), .q(
        \pipeline/regfile/data[30][24] ) );
  dp_1 \pipeline/regfile/data_reg[30][25]  ( .ip(n8943), .ck(clk), .q(
        \pipeline/regfile/data[30][25] ) );
  dp_1 \pipeline/regfile/data_reg[30][26]  ( .ip(n8942), .ck(clk), .q(
        \pipeline/regfile/data[30][26] ) );
  dp_1 \pipeline/regfile/data_reg[30][27]  ( .ip(n8941), .ck(clk), .q(
        \pipeline/regfile/data[30][27] ) );
  dp_1 \pipeline/regfile/data_reg[30][28]  ( .ip(n8940), .ck(clk), .q(
        \pipeline/regfile/data[30][28] ) );
  dp_1 \pipeline/regfile/data_reg[30][29]  ( .ip(n8939), .ck(clk), .q(
        \pipeline/regfile/data[30][29] ) );
  dp_1 \pipeline/regfile/data_reg[30][30]  ( .ip(n8938), .ck(clk), .q(
        \pipeline/regfile/data[30][30] ) );
  dp_1 \pipeline/regfile/data_reg[30][31]  ( .ip(n8937), .ck(clk), .q(
        \pipeline/regfile/data[30][31] ) );
  dp_1 \pipeline/regfile/data_reg[31][0]  ( .ip(n8936), .ck(clk), .q(
        \pipeline/regfile/data[31][0] ) );
  dp_1 \pipeline/regfile/data_reg[31][1]  ( .ip(n8935), .ck(clk), .q(
        \pipeline/regfile/data[31][1] ) );
  dp_1 \pipeline/regfile/data_reg[31][2]  ( .ip(n8934), .ck(clk), .q(
        \pipeline/regfile/data[31][2] ) );
  dp_1 \pipeline/regfile/data_reg[31][3]  ( .ip(n8933), .ck(clk), .q(
        \pipeline/regfile/data[31][3] ) );
  dp_1 \pipeline/regfile/data_reg[31][4]  ( .ip(n8932), .ck(clk), .q(
        \pipeline/regfile/data[31][4] ) );
  dp_1 \pipeline/regfile/data_reg[31][5]  ( .ip(n8931), .ck(clk), .q(
        \pipeline/regfile/data[31][5] ) );
  dp_1 \pipeline/regfile/data_reg[31][6]  ( .ip(n8930), .ck(clk), .q(
        \pipeline/regfile/data[31][6] ) );
  dp_1 \pipeline/regfile/data_reg[31][7]  ( .ip(n8929), .ck(clk), .q(
        \pipeline/regfile/data[31][7] ) );
  dp_1 \pipeline/regfile/data_reg[31][8]  ( .ip(n8928), .ck(clk), .q(
        \pipeline/regfile/data[31][8] ) );
  dp_1 \pipeline/regfile/data_reg[31][9]  ( .ip(n8927), .ck(clk), .q(
        \pipeline/regfile/data[31][9] ) );
  dp_1 \pipeline/regfile/data_reg[31][10]  ( .ip(n8926), .ck(clk), .q(
        \pipeline/regfile/data[31][10] ) );
  dp_1 \pipeline/regfile/data_reg[31][11]  ( .ip(n8925), .ck(clk), .q(
        \pipeline/regfile/data[31][11] ) );
  dp_1 \pipeline/regfile/data_reg[31][12]  ( .ip(n8924), .ck(clk), .q(
        \pipeline/regfile/data[31][12] ) );
  dp_1 \pipeline/regfile/data_reg[31][13]  ( .ip(n8923), .ck(clk), .q(
        \pipeline/regfile/data[31][13] ) );
  dp_1 \pipeline/regfile/data_reg[31][14]  ( .ip(n8922), .ck(clk), .q(
        \pipeline/regfile/data[31][14] ) );
  dp_1 \pipeline/regfile/data_reg[31][15]  ( .ip(n8921), .ck(clk), .q(
        \pipeline/regfile/data[31][15] ) );
  dp_1 \pipeline/regfile/data_reg[31][16]  ( .ip(n8920), .ck(clk), .q(
        \pipeline/regfile/data[31][16] ) );
  dp_1 \pipeline/regfile/data_reg[31][17]  ( .ip(n8919), .ck(clk), .q(
        \pipeline/regfile/data[31][17] ) );
  dp_1 \pipeline/regfile/data_reg[31][18]  ( .ip(n8918), .ck(clk), .q(
        \pipeline/regfile/data[31][18] ) );
  dp_1 \pipeline/regfile/data_reg[31][19]  ( .ip(n8917), .ck(clk), .q(
        \pipeline/regfile/data[31][19] ) );
  dp_1 \pipeline/regfile/data_reg[31][20]  ( .ip(n8916), .ck(clk), .q(
        \pipeline/regfile/data[31][20] ) );
  dp_1 \pipeline/regfile/data_reg[31][21]  ( .ip(n8915), .ck(clk), .q(
        \pipeline/regfile/data[31][21] ) );
  dp_1 \pipeline/regfile/data_reg[31][22]  ( .ip(n8914), .ck(clk), .q(
        \pipeline/regfile/data[31][22] ) );
  dp_1 \pipeline/regfile/data_reg[31][23]  ( .ip(n8913), .ck(clk), .q(
        \pipeline/regfile/data[31][23] ) );
  dp_1 \pipeline/regfile/data_reg[31][24]  ( .ip(n8912), .ck(clk), .q(
        \pipeline/regfile/data[31][24] ) );
  dp_1 \pipeline/regfile/data_reg[31][25]  ( .ip(n8911), .ck(clk), .q(
        \pipeline/regfile/data[31][25] ) );
  dp_1 \pipeline/regfile/data_reg[31][26]  ( .ip(n8910), .ck(clk), .q(
        \pipeline/regfile/data[31][26] ) );
  dp_1 \pipeline/regfile/data_reg[31][27]  ( .ip(n8909), .ck(clk), .q(
        \pipeline/regfile/data[31][27] ) );
  dp_1 \pipeline/regfile/data_reg[31][28]  ( .ip(n8908), .ck(clk), .q(
        \pipeline/regfile/data[31][28] ) );
  dp_1 \pipeline/regfile/data_reg[31][29]  ( .ip(n8907), .ck(clk), .q(
        \pipeline/regfile/data[31][29] ) );
  dp_1 \pipeline/regfile/data_reg[31][30]  ( .ip(n8906), .ck(clk), .q(
        \pipeline/regfile/data[31][30] ) );
  dp_1 \pipeline/regfile/data_reg[31][31]  ( .ip(n8905), .ck(clk), .q(
        \pipeline/regfile/data[31][31] ) );
  dp_1 \pipeline/ctrl/wb_src_sel_WB_reg[1]  ( .ip(n10065), .ck(clk), .q(
        \pipeline/wb_src_sel_WB [1]) );
  dp_1 \pipeline/ctrl/wb_src_sel_WB_reg[0]  ( .ip(n10066), .ck(clk), .q(
        \pipeline/wb_src_sel_WB [0]) );
  dp_1 \pipeline/ctrl/replay_IF_reg  ( .ip(\pipeline/ctrl/N66 ), .ck(clk), .q(
        \pipeline/ctrl/replay_IF ) );
  dp_1 \pipeline/store_data_WB_reg[31]  ( .ip(n8808), .ck(clk), .q(
        \pipeline/store_data_WB [31]) );
  dp_1 \pipeline/csr/mie_reg[0]  ( .ip(n10060), .ck(clk), .q(
        \pipeline/csr/mie [0]) );
  dp_1 \pipeline/csr/mie_reg[1]  ( .ip(n10059), .ck(clk), .q(
        \pipeline/csr/mie [1]) );
  dp_1 \pipeline/csr/mie_reg[2]  ( .ip(n10058), .ck(clk), .q(
        \pipeline/csr/mie [2]) );
  dp_1 \pipeline/csr/mie_reg[3]  ( .ip(n10057), .ck(clk), .q(
        \pipeline/csr/mie [3]) );
  dp_1 \pipeline/csr/mie_reg[4]  ( .ip(n10056), .ck(clk), .q(
        \pipeline/csr/mie [4]) );
  dp_1 \pipeline/csr/mie_reg[5]  ( .ip(n10055), .ck(clk), .q(
        \pipeline/csr/mie [5]) );
  dp_1 \pipeline/csr/mie_reg[6]  ( .ip(n10054), .ck(clk), .q(
        \pipeline/csr/mie [6]) );
  dp_1 \pipeline/csr/mie_reg[7]  ( .ip(n10053), .ck(clk), .q(
        \pipeline/csr/mie [7]) );
  dp_1 \pipeline/csr/mie_reg[8]  ( .ip(n10052), .ck(clk), .q(
        \pipeline/csr/mie [8]) );
  dp_1 \pipeline/csr/mie_reg[9]  ( .ip(n10051), .ck(clk), .q(
        \pipeline/csr/mie [9]) );
  dp_1 \pipeline/csr/mie_reg[10]  ( .ip(n10050), .ck(clk), .q(
        \pipeline/csr/mie [10]) );
  dp_1 \pipeline/csr/mie_reg[11]  ( .ip(n10049), .ck(clk), .q(
        \pipeline/csr/mie [11]) );
  dp_1 \pipeline/csr/mie_reg[12]  ( .ip(n10048), .ck(clk), .q(
        \pipeline/csr/mie [12]) );
  dp_1 \pipeline/csr/mie_reg[13]  ( .ip(n10047), .ck(clk), .q(
        \pipeline/csr/mie [13]) );
  dp_1 \pipeline/csr/mie_reg[14]  ( .ip(n10046), .ck(clk), .q(
        \pipeline/csr/mie [14]) );
  dp_1 \pipeline/csr/mie_reg[15]  ( .ip(n10045), .ck(clk), .q(
        \pipeline/csr/mie [15]) );
  dp_1 \pipeline/csr/mie_reg[16]  ( .ip(n10044), .ck(clk), .q(
        \pipeline/csr/mie [16]) );
  dp_1 \pipeline/csr/mie_reg[17]  ( .ip(n10043), .ck(clk), .q(
        \pipeline/csr/mie [17]) );
  dp_1 \pipeline/csr/mie_reg[18]  ( .ip(n10042), .ck(clk), .q(
        \pipeline/csr/mie [18]) );
  dp_1 \pipeline/csr/mie_reg[19]  ( .ip(n10041), .ck(clk), .q(
        \pipeline/csr/mie [19]) );
  dp_1 \pipeline/csr/mie_reg[20]  ( .ip(n10040), .ck(clk), .q(
        \pipeline/csr/mie [20]) );
  dp_1 \pipeline/csr/mie_reg[21]  ( .ip(n10039), .ck(clk), .q(
        \pipeline/csr/mie [21]) );
  dp_1 \pipeline/csr/mie_reg[22]  ( .ip(n10038), .ck(clk), .q(
        \pipeline/csr/mie [22]) );
  dp_1 \pipeline/csr/mie_reg[23]  ( .ip(n10037), .ck(clk), .q(
        \pipeline/csr/mie [23]) );
  dp_1 \pipeline/csr/mie_reg[24]  ( .ip(n10036), .ck(clk), .q(
        \pipeline/csr/mie [24]) );
  dp_1 \pipeline/csr/mie_reg[25]  ( .ip(n10035), .ck(clk), .q(
        \pipeline/csr/mie [25]) );
  dp_1 \pipeline/csr/mie_reg[26]  ( .ip(n10034), .ck(clk), .q(
        \pipeline/csr/mie [26]) );
  dp_1 \pipeline/csr/mie_reg[27]  ( .ip(n10033), .ck(clk), .q(
        \pipeline/csr/mie [27]) );
  dp_1 \pipeline/csr/mie_reg[28]  ( .ip(n10032), .ck(clk), .q(
        \pipeline/csr/mie [28]) );
  dp_1 \pipeline/csr/mie_reg[29]  ( .ip(n10031), .ck(clk), .q(
        \pipeline/csr/mie [29]) );
  dp_1 \pipeline/csr/mie_reg[30]  ( .ip(n10030), .ck(clk), .q(
        \pipeline/csr/mie [30]) );
  dp_1 \pipeline/csr/mie_reg[31]  ( .ip(n10029), .ck(clk), .q(
        \pipeline/csr/mie [31]) );
  dp_1 \pipeline/csr/mtime_full_reg[0]  ( .ip(\pipeline/csr/N2081 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [0]) );
  dp_1 \pipeline/csr/mtime_full_reg[1]  ( .ip(\pipeline/csr/N2082 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [1]) );
  dp_1 \pipeline/csr/mtime_full_reg[2]  ( .ip(\pipeline/csr/N2083 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [2]) );
  dp_1 \pipeline/csr/mtime_full_reg[3]  ( .ip(\pipeline/csr/N2084 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [3]) );
  dp_1 \pipeline/csr/mtime_full_reg[4]  ( .ip(\pipeline/csr/N2085 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [4]) );
  dp_1 \pipeline/csr/mtime_full_reg[5]  ( .ip(\pipeline/csr/N2086 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [5]) );
  dp_1 \pipeline/csr/mtime_full_reg[6]  ( .ip(\pipeline/csr/N2087 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [6]) );
  dp_1 \pipeline/csr/mtime_full_reg[7]  ( .ip(\pipeline/csr/N2088 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [7]) );
  dp_1 \pipeline/csr/mtime_full_reg[8]  ( .ip(\pipeline/csr/N2089 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [8]) );
  dp_1 \pipeline/csr/mtime_full_reg[9]  ( .ip(\pipeline/csr/N2090 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [9]) );
  dp_1 \pipeline/csr/mtime_full_reg[10]  ( .ip(\pipeline/csr/N2091 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [10]) );
  dp_1 \pipeline/csr/mtime_full_reg[11]  ( .ip(\pipeline/csr/N2092 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [11]) );
  dp_1 \pipeline/csr/mtime_full_reg[12]  ( .ip(\pipeline/csr/N2093 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [12]) );
  dp_1 \pipeline/csr/mtime_full_reg[13]  ( .ip(\pipeline/csr/N2094 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [13]) );
  dp_1 \pipeline/csr/mtime_full_reg[14]  ( .ip(\pipeline/csr/N2095 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [14]) );
  dp_1 \pipeline/csr/mtime_full_reg[15]  ( .ip(\pipeline/csr/N2096 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [15]) );
  dp_1 \pipeline/csr/mtime_full_reg[16]  ( .ip(\pipeline/csr/N2097 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [16]) );
  dp_1 \pipeline/csr/mtime_full_reg[17]  ( .ip(\pipeline/csr/N2098 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [17]) );
  dp_1 \pipeline/csr/mtime_full_reg[18]  ( .ip(\pipeline/csr/N2099 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [18]) );
  dp_1 \pipeline/csr/mtime_full_reg[19]  ( .ip(\pipeline/csr/N2100 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [19]) );
  dp_1 \pipeline/csr/mtime_full_reg[20]  ( .ip(\pipeline/csr/N2101 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [20]) );
  dp_1 \pipeline/csr/mtime_full_reg[21]  ( .ip(\pipeline/csr/N2102 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [21]) );
  dp_1 \pipeline/csr/mtime_full_reg[22]  ( .ip(\pipeline/csr/N2103 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [22]) );
  dp_1 \pipeline/csr/mtime_full_reg[23]  ( .ip(\pipeline/csr/N2104 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [23]) );
  dp_1 \pipeline/csr/mtime_full_reg[24]  ( .ip(\pipeline/csr/N2105 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [24]) );
  dp_1 \pipeline/csr/mtime_full_reg[25]  ( .ip(\pipeline/csr/N2106 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [25]) );
  dp_1 \pipeline/csr/mtime_full_reg[26]  ( .ip(\pipeline/csr/N2107 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [26]) );
  dp_1 \pipeline/csr/mtime_full_reg[27]  ( .ip(\pipeline/csr/N2108 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [27]) );
  dp_1 \pipeline/csr/mtime_full_reg[28]  ( .ip(\pipeline/csr/N2109 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [28]) );
  dp_1 \pipeline/csr/mtime_full_reg[29]  ( .ip(\pipeline/csr/N2110 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [29]) );
  dp_1 \pipeline/csr/mtime_full_reg[30]  ( .ip(\pipeline/csr/N2111 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [30]) );
  dp_1 \pipeline/csr/mtime_full_reg[31]  ( .ip(\pipeline/csr/N2112 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [31]) );
  dp_1 \pipeline/csr/mtime_full_reg[32]  ( .ip(\pipeline/csr/N2113 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [32]) );
  dp_1 \pipeline/csr/mtime_full_reg[33]  ( .ip(\pipeline/csr/N2114 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [33]) );
  dp_1 \pipeline/csr/mtime_full_reg[34]  ( .ip(\pipeline/csr/N2115 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [34]) );
  dp_1 \pipeline/csr/mtime_full_reg[35]  ( .ip(\pipeline/csr/N2116 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [35]) );
  dp_1 \pipeline/csr/mtime_full_reg[36]  ( .ip(\pipeline/csr/N2117 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [36]) );
  dp_1 \pipeline/csr/mtime_full_reg[37]  ( .ip(\pipeline/csr/N2118 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [37]) );
  dp_1 \pipeline/csr/mtime_full_reg[38]  ( .ip(\pipeline/csr/N2119 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [38]) );
  dp_1 \pipeline/csr/mtime_full_reg[39]  ( .ip(\pipeline/csr/N2120 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [39]) );
  dp_1 \pipeline/csr/mtime_full_reg[40]  ( .ip(\pipeline/csr/N2121 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [40]) );
  dp_1 \pipeline/csr/mtime_full_reg[41]  ( .ip(\pipeline/csr/N2122 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [41]) );
  dp_1 \pipeline/csr/mtime_full_reg[42]  ( .ip(\pipeline/csr/N2123 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [42]) );
  dp_1 \pipeline/csr/mtime_full_reg[43]  ( .ip(\pipeline/csr/N2124 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [43]) );
  dp_1 \pipeline/csr/mtime_full_reg[44]  ( .ip(\pipeline/csr/N2125 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [44]) );
  dp_1 \pipeline/csr/mtime_full_reg[45]  ( .ip(\pipeline/csr/N2126 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [45]) );
  dp_1 \pipeline/csr/mtime_full_reg[46]  ( .ip(\pipeline/csr/N2127 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [46]) );
  dp_1 \pipeline/csr/mtime_full_reg[47]  ( .ip(\pipeline/csr/N2128 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [47]) );
  dp_1 \pipeline/csr/mtime_full_reg[48]  ( .ip(\pipeline/csr/N2129 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [48]) );
  dp_1 \pipeline/csr/mtime_full_reg[49]  ( .ip(\pipeline/csr/N2130 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [49]) );
  dp_1 \pipeline/csr/mtime_full_reg[50]  ( .ip(\pipeline/csr/N2131 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [50]) );
  dp_1 \pipeline/csr/mtime_full_reg[51]  ( .ip(\pipeline/csr/N2132 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [51]) );
  dp_1 \pipeline/csr/mtime_full_reg[52]  ( .ip(\pipeline/csr/N2133 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [52]) );
  dp_1 \pipeline/csr/mtime_full_reg[53]  ( .ip(\pipeline/csr/N2134 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [53]) );
  dp_1 \pipeline/csr/mtime_full_reg[54]  ( .ip(\pipeline/csr/N2135 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [54]) );
  dp_1 \pipeline/csr/mtime_full_reg[55]  ( .ip(\pipeline/csr/N2136 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [55]) );
  dp_1 \pipeline/csr/mtime_full_reg[56]  ( .ip(\pipeline/csr/N2137 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [56]) );
  dp_1 \pipeline/csr/mtime_full_reg[57]  ( .ip(\pipeline/csr/N2138 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [57]) );
  dp_1 \pipeline/csr/mtime_full_reg[58]  ( .ip(\pipeline/csr/N2139 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [58]) );
  dp_1 \pipeline/csr/mtime_full_reg[59]  ( .ip(\pipeline/csr/N2140 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [59]) );
  dp_1 \pipeline/csr/mtime_full_reg[60]  ( .ip(\pipeline/csr/N2141 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [60]) );
  dp_1 \pipeline/csr/mtime_full_reg[61]  ( .ip(\pipeline/csr/N2142 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [61]) );
  dp_1 \pipeline/csr/mtime_full_reg[62]  ( .ip(\pipeline/csr/N2143 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [62]) );
  dp_1 \pipeline/csr/mtime_full_reg[63]  ( .ip(\pipeline/csr/N2144 ), .ck(clk), 
        .q(\pipeline/csr/mtime_full [63]) );
  dp_1 \pipeline/csr/time_full_reg[0]  ( .ip(\pipeline/csr/N1937 ), .ck(clk), 
        .q(\pipeline/csr/time_full [0]) );
  dp_1 \pipeline/csr/time_full_reg[1]  ( .ip(\pipeline/csr/N1938 ), .ck(clk), 
        .q(\pipeline/csr/time_full [1]) );
  dp_1 \pipeline/csr/time_full_reg[2]  ( .ip(\pipeline/csr/N1939 ), .ck(clk), 
        .q(\pipeline/csr/time_full [2]) );
  dp_1 \pipeline/csr/time_full_reg[3]  ( .ip(\pipeline/csr/N1940 ), .ck(clk), 
        .q(\pipeline/csr/time_full [3]) );
  dp_1 \pipeline/csr/time_full_reg[4]  ( .ip(\pipeline/csr/N1941 ), .ck(clk), 
        .q(\pipeline/csr/time_full [4]) );
  dp_1 \pipeline/csr/time_full_reg[5]  ( .ip(\pipeline/csr/N1942 ), .ck(clk), 
        .q(\pipeline/csr/time_full [5]) );
  dp_1 \pipeline/csr/time_full_reg[6]  ( .ip(\pipeline/csr/N1943 ), .ck(clk), 
        .q(\pipeline/csr/time_full [6]) );
  dp_1 \pipeline/csr/time_full_reg[7]  ( .ip(\pipeline/csr/N1944 ), .ck(clk), 
        .q(\pipeline/csr/time_full [7]) );
  dp_1 \pipeline/csr/time_full_reg[8]  ( .ip(\pipeline/csr/N1945 ), .ck(clk), 
        .q(\pipeline/csr/time_full [8]) );
  dp_1 \pipeline/csr/time_full_reg[9]  ( .ip(\pipeline/csr/N1946 ), .ck(clk), 
        .q(\pipeline/csr/time_full [9]) );
  dp_1 \pipeline/csr/time_full_reg[10]  ( .ip(\pipeline/csr/N1947 ), .ck(clk), 
        .q(\pipeline/csr/time_full [10]) );
  dp_1 \pipeline/csr/time_full_reg[11]  ( .ip(\pipeline/csr/N1948 ), .ck(clk), 
        .q(\pipeline/csr/time_full [11]) );
  dp_1 \pipeline/csr/time_full_reg[12]  ( .ip(\pipeline/csr/N1949 ), .ck(clk), 
        .q(\pipeline/csr/time_full [12]) );
  dp_1 \pipeline/csr/time_full_reg[13]  ( .ip(\pipeline/csr/N1950 ), .ck(clk), 
        .q(\pipeline/csr/time_full [13]) );
  dp_1 \pipeline/csr/time_full_reg[14]  ( .ip(\pipeline/csr/N1951 ), .ck(clk), 
        .q(\pipeline/csr/time_full [14]) );
  dp_1 \pipeline/csr/time_full_reg[15]  ( .ip(\pipeline/csr/N1952 ), .ck(clk), 
        .q(\pipeline/csr/time_full [15]) );
  dp_1 \pipeline/csr/time_full_reg[16]  ( .ip(\pipeline/csr/N1953 ), .ck(clk), 
        .q(\pipeline/csr/time_full [16]) );
  dp_1 \pipeline/csr/time_full_reg[17]  ( .ip(\pipeline/csr/N1954 ), .ck(clk), 
        .q(\pipeline/csr/time_full [17]) );
  dp_1 \pipeline/csr/time_full_reg[18]  ( .ip(\pipeline/csr/N1955 ), .ck(clk), 
        .q(\pipeline/csr/time_full [18]) );
  dp_1 \pipeline/csr/time_full_reg[19]  ( .ip(\pipeline/csr/N1956 ), .ck(clk), 
        .q(\pipeline/csr/time_full [19]) );
  dp_1 \pipeline/csr/time_full_reg[20]  ( .ip(\pipeline/csr/N1957 ), .ck(clk), 
        .q(\pipeline/csr/time_full [20]) );
  dp_1 \pipeline/csr/time_full_reg[21]  ( .ip(\pipeline/csr/N1958 ), .ck(clk), 
        .q(\pipeline/csr/time_full [21]) );
  dp_1 \pipeline/csr/time_full_reg[22]  ( .ip(\pipeline/csr/N1959 ), .ck(clk), 
        .q(\pipeline/csr/time_full [22]) );
  dp_1 \pipeline/csr/time_full_reg[23]  ( .ip(\pipeline/csr/N1960 ), .ck(clk), 
        .q(\pipeline/csr/time_full [23]) );
  dp_1 \pipeline/csr/time_full_reg[24]  ( .ip(\pipeline/csr/N1961 ), .ck(clk), 
        .q(\pipeline/csr/time_full [24]) );
  dp_1 \pipeline/csr/time_full_reg[25]  ( .ip(\pipeline/csr/N1962 ), .ck(clk), 
        .q(\pipeline/csr/time_full [25]) );
  dp_1 \pipeline/csr/time_full_reg[26]  ( .ip(\pipeline/csr/N1963 ), .ck(clk), 
        .q(\pipeline/csr/time_full [26]) );
  dp_1 \pipeline/csr/time_full_reg[27]  ( .ip(\pipeline/csr/N1964 ), .ck(clk), 
        .q(\pipeline/csr/time_full [27]) );
  dp_1 \pipeline/csr/time_full_reg[28]  ( .ip(\pipeline/csr/N1965 ), .ck(clk), 
        .q(\pipeline/csr/time_full [28]) );
  dp_1 \pipeline/csr/time_full_reg[29]  ( .ip(\pipeline/csr/N1966 ), .ck(clk), 
        .q(\pipeline/csr/time_full [29]) );
  dp_1 \pipeline/csr/time_full_reg[30]  ( .ip(\pipeline/csr/N1967 ), .ck(clk), 
        .q(\pipeline/csr/time_full [30]) );
  dp_1 \pipeline/csr/time_full_reg[31]  ( .ip(\pipeline/csr/N1968 ), .ck(clk), 
        .q(\pipeline/csr/time_full [31]) );
  dp_1 \pipeline/csr/time_full_reg[32]  ( .ip(\pipeline/csr/N1969 ), .ck(clk), 
        .q(\pipeline/csr/time_full [32]) );
  dp_1 \pipeline/csr/time_full_reg[33]  ( .ip(\pipeline/csr/N1970 ), .ck(clk), 
        .q(\pipeline/csr/time_full [33]) );
  dp_1 \pipeline/csr/time_full_reg[34]  ( .ip(\pipeline/csr/N1971 ), .ck(clk), 
        .q(\pipeline/csr/time_full [34]) );
  dp_1 \pipeline/csr/time_full_reg[35]  ( .ip(\pipeline/csr/N1972 ), .ck(clk), 
        .q(\pipeline/csr/time_full [35]) );
  dp_1 \pipeline/csr/time_full_reg[36]  ( .ip(\pipeline/csr/N1973 ), .ck(clk), 
        .q(\pipeline/csr/time_full [36]) );
  dp_1 \pipeline/csr/time_full_reg[37]  ( .ip(\pipeline/csr/N1974 ), .ck(clk), 
        .q(\pipeline/csr/time_full [37]) );
  dp_1 \pipeline/csr/time_full_reg[38]  ( .ip(\pipeline/csr/N1975 ), .ck(clk), 
        .q(\pipeline/csr/time_full [38]) );
  dp_1 \pipeline/csr/time_full_reg[39]  ( .ip(\pipeline/csr/N1976 ), .ck(clk), 
        .q(\pipeline/csr/time_full [39]) );
  dp_1 \pipeline/csr/time_full_reg[40]  ( .ip(\pipeline/csr/N1977 ), .ck(clk), 
        .q(\pipeline/csr/time_full [40]) );
  dp_1 \pipeline/csr/time_full_reg[41]  ( .ip(\pipeline/csr/N1978 ), .ck(clk), 
        .q(\pipeline/csr/time_full [41]) );
  dp_1 \pipeline/csr/time_full_reg[42]  ( .ip(\pipeline/csr/N1979 ), .ck(clk), 
        .q(\pipeline/csr/time_full [42]) );
  dp_1 \pipeline/csr/time_full_reg[43]  ( .ip(\pipeline/csr/N1980 ), .ck(clk), 
        .q(\pipeline/csr/time_full [43]) );
  dp_1 \pipeline/csr/time_full_reg[44]  ( .ip(\pipeline/csr/N1981 ), .ck(clk), 
        .q(\pipeline/csr/time_full [44]) );
  dp_1 \pipeline/csr/time_full_reg[45]  ( .ip(\pipeline/csr/N1982 ), .ck(clk), 
        .q(\pipeline/csr/time_full [45]) );
  dp_1 \pipeline/csr/time_full_reg[46]  ( .ip(\pipeline/csr/N1983 ), .ck(clk), 
        .q(\pipeline/csr/time_full [46]) );
  dp_1 \pipeline/csr/time_full_reg[47]  ( .ip(\pipeline/csr/N1984 ), .ck(clk), 
        .q(\pipeline/csr/time_full [47]) );
  dp_1 \pipeline/csr/time_full_reg[48]  ( .ip(\pipeline/csr/N1985 ), .ck(clk), 
        .q(\pipeline/csr/time_full [48]) );
  dp_1 \pipeline/csr/time_full_reg[49]  ( .ip(\pipeline/csr/N1986 ), .ck(clk), 
        .q(\pipeline/csr/time_full [49]) );
  dp_1 \pipeline/csr/time_full_reg[50]  ( .ip(\pipeline/csr/N1987 ), .ck(clk), 
        .q(\pipeline/csr/time_full [50]) );
  dp_1 \pipeline/csr/time_full_reg[51]  ( .ip(\pipeline/csr/N1988 ), .ck(clk), 
        .q(\pipeline/csr/time_full [51]) );
  dp_1 \pipeline/csr/time_full_reg[52]  ( .ip(\pipeline/csr/N1989 ), .ck(clk), 
        .q(\pipeline/csr/time_full [52]) );
  dp_1 \pipeline/csr/time_full_reg[53]  ( .ip(\pipeline/csr/N1990 ), .ck(clk), 
        .q(\pipeline/csr/time_full [53]) );
  dp_1 \pipeline/csr/time_full_reg[54]  ( .ip(\pipeline/csr/N1991 ), .ck(clk), 
        .q(\pipeline/csr/time_full [54]) );
  dp_1 \pipeline/csr/time_full_reg[55]  ( .ip(\pipeline/csr/N1992 ), .ck(clk), 
        .q(\pipeline/csr/time_full [55]) );
  dp_1 \pipeline/csr/time_full_reg[56]  ( .ip(\pipeline/csr/N1993 ), .ck(clk), 
        .q(\pipeline/csr/time_full [56]) );
  dp_1 \pipeline/csr/time_full_reg[57]  ( .ip(\pipeline/csr/N1994 ), .ck(clk), 
        .q(\pipeline/csr/time_full [57]) );
  dp_1 \pipeline/csr/time_full_reg[58]  ( .ip(\pipeline/csr/N1995 ), .ck(clk), 
        .q(\pipeline/csr/time_full [58]) );
  dp_1 \pipeline/csr/time_full_reg[59]  ( .ip(\pipeline/csr/N1996 ), .ck(clk), 
        .q(\pipeline/csr/time_full [59]) );
  dp_1 \pipeline/csr/time_full_reg[60]  ( .ip(\pipeline/csr/N1997 ), .ck(clk), 
        .q(\pipeline/csr/time_full [60]) );
  dp_1 \pipeline/csr/time_full_reg[61]  ( .ip(\pipeline/csr/N1998 ), .ck(clk), 
        .q(\pipeline/csr/time_full [61]) );
  dp_1 \pipeline/csr/time_full_reg[62]  ( .ip(\pipeline/csr/N1999 ), .ck(clk), 
        .q(\pipeline/csr/time_full [62]) );
  dp_1 \pipeline/csr/time_full_reg[63]  ( .ip(\pipeline/csr/N2000 ), .ck(clk), 
        .q(\pipeline/csr/time_full [63]) );
  dp_1 \pipeline/csr/cycle_full_reg[0]  ( .ip(\pipeline/csr/N1873 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [0]) );
  dp_1 \pipeline/csr/cycle_full_reg[1]  ( .ip(\pipeline/csr/N1874 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [1]) );
  dp_1 \pipeline/csr/cycle_full_reg[2]  ( .ip(\pipeline/csr/N1875 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [2]) );
  dp_1 \pipeline/csr/cycle_full_reg[3]  ( .ip(\pipeline/csr/N1876 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [3]) );
  dp_1 \pipeline/csr/cycle_full_reg[4]  ( .ip(\pipeline/csr/N1877 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [4]) );
  dp_1 \pipeline/csr/cycle_full_reg[5]  ( .ip(\pipeline/csr/N1878 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [5]) );
  dp_1 \pipeline/csr/cycle_full_reg[6]  ( .ip(\pipeline/csr/N1879 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [6]) );
  dp_1 \pipeline/csr/cycle_full_reg[7]  ( .ip(\pipeline/csr/N1880 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [7]) );
  dp_1 \pipeline/csr/cycle_full_reg[8]  ( .ip(\pipeline/csr/N1881 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [8]) );
  dp_1 \pipeline/csr/cycle_full_reg[9]  ( .ip(\pipeline/csr/N1882 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [9]) );
  dp_1 \pipeline/csr/cycle_full_reg[10]  ( .ip(\pipeline/csr/N1883 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [10]) );
  dp_1 \pipeline/csr/cycle_full_reg[11]  ( .ip(\pipeline/csr/N1884 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [11]) );
  dp_1 \pipeline/csr/cycle_full_reg[12]  ( .ip(\pipeline/csr/N1885 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [12]) );
  dp_1 \pipeline/csr/cycle_full_reg[13]  ( .ip(\pipeline/csr/N1886 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [13]) );
  dp_1 \pipeline/csr/cycle_full_reg[14]  ( .ip(\pipeline/csr/N1887 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [14]) );
  dp_1 \pipeline/csr/cycle_full_reg[15]  ( .ip(\pipeline/csr/N1888 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [15]) );
  dp_1 \pipeline/csr/cycle_full_reg[16]  ( .ip(\pipeline/csr/N1889 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [16]) );
  dp_1 \pipeline/csr/cycle_full_reg[17]  ( .ip(\pipeline/csr/N1890 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [17]) );
  dp_1 \pipeline/csr/cycle_full_reg[18]  ( .ip(\pipeline/csr/N1891 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [18]) );
  dp_1 \pipeline/csr/cycle_full_reg[19]  ( .ip(\pipeline/csr/N1892 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [19]) );
  dp_1 \pipeline/csr/cycle_full_reg[20]  ( .ip(\pipeline/csr/N1893 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [20]) );
  dp_1 \pipeline/csr/cycle_full_reg[21]  ( .ip(\pipeline/csr/N1894 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [21]) );
  dp_1 \pipeline/csr/cycle_full_reg[22]  ( .ip(\pipeline/csr/N1895 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [22]) );
  dp_1 \pipeline/csr/cycle_full_reg[23]  ( .ip(\pipeline/csr/N1896 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [23]) );
  dp_1 \pipeline/csr/cycle_full_reg[24]  ( .ip(\pipeline/csr/N1897 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [24]) );
  dp_1 \pipeline/csr/cycle_full_reg[25]  ( .ip(\pipeline/csr/N1898 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [25]) );
  dp_1 \pipeline/csr/cycle_full_reg[26]  ( .ip(\pipeline/csr/N1899 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [26]) );
  dp_1 \pipeline/csr/cycle_full_reg[27]  ( .ip(\pipeline/csr/N1900 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [27]) );
  dp_1 \pipeline/csr/cycle_full_reg[28]  ( .ip(\pipeline/csr/N1901 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [28]) );
  dp_1 \pipeline/csr/cycle_full_reg[29]  ( .ip(\pipeline/csr/N1902 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [29]) );
  dp_1 \pipeline/csr/cycle_full_reg[30]  ( .ip(\pipeline/csr/N1903 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [30]) );
  dp_1 \pipeline/csr/cycle_full_reg[31]  ( .ip(\pipeline/csr/N1904 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [31]) );
  dp_1 \pipeline/csr/cycle_full_reg[32]  ( .ip(\pipeline/csr/N1905 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [32]) );
  dp_1 \pipeline/csr/cycle_full_reg[33]  ( .ip(\pipeline/csr/N1906 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [33]) );
  dp_1 \pipeline/csr/cycle_full_reg[34]  ( .ip(\pipeline/csr/N1907 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [34]) );
  dp_1 \pipeline/csr/cycle_full_reg[35]  ( .ip(\pipeline/csr/N1908 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [35]) );
  dp_1 \pipeline/csr/cycle_full_reg[36]  ( .ip(\pipeline/csr/N1909 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [36]) );
  dp_1 \pipeline/csr/cycle_full_reg[37]  ( .ip(\pipeline/csr/N1910 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [37]) );
  dp_1 \pipeline/csr/cycle_full_reg[38]  ( .ip(\pipeline/csr/N1911 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [38]) );
  dp_1 \pipeline/csr/cycle_full_reg[39]  ( .ip(\pipeline/csr/N1912 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [39]) );
  dp_1 \pipeline/csr/cycle_full_reg[40]  ( .ip(\pipeline/csr/N1913 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [40]) );
  dp_1 \pipeline/csr/cycle_full_reg[41]  ( .ip(\pipeline/csr/N1914 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [41]) );
  dp_1 \pipeline/csr/cycle_full_reg[42]  ( .ip(\pipeline/csr/N1915 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [42]) );
  dp_1 \pipeline/csr/cycle_full_reg[43]  ( .ip(\pipeline/csr/N1916 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [43]) );
  dp_1 \pipeline/csr/cycle_full_reg[44]  ( .ip(\pipeline/csr/N1917 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [44]) );
  dp_1 \pipeline/csr/cycle_full_reg[45]  ( .ip(\pipeline/csr/N1918 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [45]) );
  dp_1 \pipeline/csr/cycle_full_reg[46]  ( .ip(\pipeline/csr/N1919 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [46]) );
  dp_1 \pipeline/csr/cycle_full_reg[47]  ( .ip(\pipeline/csr/N1920 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [47]) );
  dp_1 \pipeline/csr/cycle_full_reg[48]  ( .ip(\pipeline/csr/N1921 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [48]) );
  dp_1 \pipeline/csr/cycle_full_reg[49]  ( .ip(\pipeline/csr/N1922 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [49]) );
  dp_1 \pipeline/csr/cycle_full_reg[50]  ( .ip(\pipeline/csr/N1923 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [50]) );
  dp_1 \pipeline/csr/cycle_full_reg[51]  ( .ip(\pipeline/csr/N1924 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [51]) );
  dp_1 \pipeline/csr/cycle_full_reg[52]  ( .ip(\pipeline/csr/N1925 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [52]) );
  dp_1 \pipeline/csr/cycle_full_reg[53]  ( .ip(\pipeline/csr/N1926 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [53]) );
  dp_1 \pipeline/csr/cycle_full_reg[54]  ( .ip(\pipeline/csr/N1927 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [54]) );
  dp_1 \pipeline/csr/cycle_full_reg[55]  ( .ip(\pipeline/csr/N1928 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [55]) );
  dp_1 \pipeline/csr/cycle_full_reg[56]  ( .ip(\pipeline/csr/N1929 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [56]) );
  dp_1 \pipeline/csr/cycle_full_reg[57]  ( .ip(\pipeline/csr/N1930 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [57]) );
  dp_1 \pipeline/csr/cycle_full_reg[58]  ( .ip(\pipeline/csr/N1931 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [58]) );
  dp_1 \pipeline/csr/cycle_full_reg[59]  ( .ip(\pipeline/csr/N1932 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [59]) );
  dp_1 \pipeline/csr/cycle_full_reg[60]  ( .ip(\pipeline/csr/N1933 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [60]) );
  dp_1 \pipeline/csr/cycle_full_reg[61]  ( .ip(\pipeline/csr/N1934 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [61]) );
  dp_1 \pipeline/csr/cycle_full_reg[62]  ( .ip(\pipeline/csr/N1935 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [62]) );
  dp_1 \pipeline/csr/cycle_full_reg[63]  ( .ip(\pipeline/csr/N1936 ), .ck(clk), 
        .q(\pipeline/csr/cycle_full [63]) );
  dp_1 \pipeline/csr/mtimecmp_reg[0]  ( .ip(n10022), .ck(clk), .q(
        \pipeline/csr/mtimecmp [0]) );
  dp_1 \pipeline/csr/mtimecmp_reg[1]  ( .ip(n10021), .ck(clk), .q(
        \pipeline/csr/mtimecmp [1]) );
  dp_1 \pipeline/csr/mtimecmp_reg[2]  ( .ip(n10020), .ck(clk), .q(
        \pipeline/csr/mtimecmp [2]) );
  dp_1 \pipeline/csr/mtimecmp_reg[3]  ( .ip(n10019), .ck(clk), .q(
        \pipeline/csr/mtimecmp [3]) );
  dp_1 \pipeline/csr/mtimecmp_reg[4]  ( .ip(n10018), .ck(clk), .q(
        \pipeline/csr/mtimecmp [4]) );
  dp_1 \pipeline/csr/mtimecmp_reg[5]  ( .ip(n10017), .ck(clk), .q(
        \pipeline/csr/mtimecmp [5]) );
  dp_1 \pipeline/csr/mtimecmp_reg[6]  ( .ip(n10016), .ck(clk), .q(
        \pipeline/csr/mtimecmp [6]) );
  dp_1 \pipeline/csr/mtimecmp_reg[7]  ( .ip(n10015), .ck(clk), .q(
        \pipeline/csr/mtimecmp [7]) );
  dp_1 \pipeline/csr/mtimecmp_reg[8]  ( .ip(n10014), .ck(clk), .q(
        \pipeline/csr/mtimecmp [8]) );
  dp_1 \pipeline/csr/mtimecmp_reg[9]  ( .ip(n10013), .ck(clk), .q(
        \pipeline/csr/mtimecmp [9]) );
  dp_1 \pipeline/csr/mtimecmp_reg[10]  ( .ip(n10012), .ck(clk), .q(
        \pipeline/csr/mtimecmp [10]) );
  dp_1 \pipeline/csr/mtimecmp_reg[11]  ( .ip(n10011), .ck(clk), .q(
        \pipeline/csr/mtimecmp [11]) );
  dp_1 \pipeline/csr/mtimecmp_reg[12]  ( .ip(n10010), .ck(clk), .q(
        \pipeline/csr/mtimecmp [12]) );
  dp_1 \pipeline/csr/mtimecmp_reg[13]  ( .ip(n10009), .ck(clk), .q(
        \pipeline/csr/mtimecmp [13]) );
  dp_1 \pipeline/csr/mtimecmp_reg[14]  ( .ip(n10008), .ck(clk), .q(
        \pipeline/csr/mtimecmp [14]) );
  dp_1 \pipeline/csr/mtimecmp_reg[15]  ( .ip(n10007), .ck(clk), .q(
        \pipeline/csr/mtimecmp [15]) );
  dp_1 \pipeline/csr/mtimecmp_reg[16]  ( .ip(n10006), .ck(clk), .q(
        \pipeline/csr/mtimecmp [16]) );
  dp_1 \pipeline/csr/mtimecmp_reg[17]  ( .ip(n10005), .ck(clk), .q(
        \pipeline/csr/mtimecmp [17]) );
  dp_1 \pipeline/csr/mtimecmp_reg[18]  ( .ip(n10004), .ck(clk), .q(
        \pipeline/csr/mtimecmp [18]) );
  dp_1 \pipeline/csr/mtimecmp_reg[19]  ( .ip(n10003), .ck(clk), .q(
        \pipeline/csr/mtimecmp [19]) );
  dp_1 \pipeline/csr/mtimecmp_reg[20]  ( .ip(n10002), .ck(clk), .q(
        \pipeline/csr/mtimecmp [20]) );
  dp_1 \pipeline/csr/mtimecmp_reg[21]  ( .ip(n10001), .ck(clk), .q(
        \pipeline/csr/mtimecmp [21]) );
  dp_1 \pipeline/csr/mtimecmp_reg[22]  ( .ip(n10000), .ck(clk), .q(
        \pipeline/csr/mtimecmp [22]) );
  dp_1 \pipeline/csr/mtimecmp_reg[23]  ( .ip(n9999), .ck(clk), .q(
        \pipeline/csr/mtimecmp [23]) );
  dp_1 \pipeline/csr/mtimecmp_reg[24]  ( .ip(n9998), .ck(clk), .q(
        \pipeline/csr/mtimecmp [24]) );
  dp_1 \pipeline/csr/mtimecmp_reg[25]  ( .ip(n9997), .ck(clk), .q(
        \pipeline/csr/mtimecmp [25]) );
  dp_1 \pipeline/csr/mtimecmp_reg[26]  ( .ip(n9996), .ck(clk), .q(
        \pipeline/csr/mtimecmp [26]) );
  dp_1 \pipeline/csr/mtimecmp_reg[27]  ( .ip(n9995), .ck(clk), .q(
        \pipeline/csr/mtimecmp [27]) );
  dp_1 \pipeline/csr/mtimecmp_reg[28]  ( .ip(n9994), .ck(clk), .q(
        \pipeline/csr/mtimecmp [28]) );
  dp_1 \pipeline/csr/mtimecmp_reg[29]  ( .ip(n9993), .ck(clk), .q(
        \pipeline/csr/mtimecmp [29]) );
  dp_1 \pipeline/csr/mtimecmp_reg[30]  ( .ip(n9992), .ck(clk), .q(
        \pipeline/csr/mtimecmp [30]) );
  dp_1 \pipeline/csr/mtimecmp_reg[31]  ( .ip(n9991), .ck(clk), .q(
        \pipeline/csr/mtimecmp [31]) );
  dp_1 \pipeline/csr/mtvec_reg[8]  ( .ip(n22857), .ck(clk), .q(
        \pipeline/csr/mtvec [8]) );
  dp_1 \pipeline/csr/mtvec_reg[2]  ( .ip(n9990), .ck(clk), .q(
        \pipeline/csr/mtvec [2]) );
  dp_1 \pipeline/csr/mtvec_reg[3]  ( .ip(n9989), .ck(clk), .q(
        \pipeline/csr/mtvec [3]) );
  dp_1 \pipeline/csr/mtvec_reg[4]  ( .ip(n9988), .ck(clk), .q(
        \pipeline/csr/mtvec [4]) );
  dp_1 \pipeline/csr/mtvec_reg[5]  ( .ip(n9987), .ck(clk), .q(
        \pipeline/csr/mtvec [5]) );
  dp_1 \pipeline/csr/mtvec_reg[6]  ( .ip(n9986), .ck(clk), .q(
        \pipeline/csr/mtvec [6]) );
  dp_1 \pipeline/csr/mtvec_reg[7]  ( .ip(n9985), .ck(clk), .q(
        \pipeline/csr/mtvec [7]) );
  dp_1 \pipeline/csr/mtvec_reg[9]  ( .ip(n9983), .ck(clk), .q(
        \pipeline/csr/mtvec [9]) );
  dp_1 \pipeline/csr/mtvec_reg[10]  ( .ip(n9982), .ck(clk), .q(
        \pipeline/csr/mtvec [10]) );
  dp_1 \pipeline/csr/mtvec_reg[11]  ( .ip(n9981), .ck(clk), .q(
        \pipeline/csr/mtvec [11]) );
  dp_1 \pipeline/csr/mtvec_reg[12]  ( .ip(n9980), .ck(clk), .q(
        \pipeline/csr/mtvec [12]) );
  dp_1 \pipeline/csr/mtvec_reg[13]  ( .ip(n9979), .ck(clk), .q(
        \pipeline/csr/mtvec [13]) );
  dp_1 \pipeline/csr/mtvec_reg[14]  ( .ip(n9978), .ck(clk), .q(
        \pipeline/csr/mtvec [14]) );
  dp_1 \pipeline/csr/mtvec_reg[15]  ( .ip(n9977), .ck(clk), .q(
        \pipeline/csr/mtvec [15]) );
  dp_1 \pipeline/csr/mtvec_reg[16]  ( .ip(n9976), .ck(clk), .q(
        \pipeline/csr/mtvec [16]) );
  dp_1 \pipeline/csr/mtvec_reg[17]  ( .ip(n9975), .ck(clk), .q(
        \pipeline/csr/mtvec [17]) );
  dp_1 \pipeline/csr/mtvec_reg[18]  ( .ip(n9974), .ck(clk), .q(
        \pipeline/csr/mtvec [18]) );
  dp_1 \pipeline/csr/mtvec_reg[19]  ( .ip(n9973), .ck(clk), .q(
        \pipeline/csr/mtvec [19]) );
  dp_1 \pipeline/csr/mtvec_reg[20]  ( .ip(n9972), .ck(clk), .q(
        \pipeline/csr/mtvec [20]) );
  dp_1 \pipeline/csr/mtvec_reg[21]  ( .ip(n9971), .ck(clk), .q(
        \pipeline/csr/mtvec [21]) );
  dp_1 \pipeline/csr/mtvec_reg[22]  ( .ip(n9970), .ck(clk), .q(
        \pipeline/csr/mtvec [22]) );
  dp_1 \pipeline/csr/mtvec_reg[23]  ( .ip(n9969), .ck(clk), .q(
        \pipeline/csr/mtvec [23]) );
  dp_1 \pipeline/csr/mtvec_reg[24]  ( .ip(n9968), .ck(clk), .q(
        \pipeline/csr/mtvec [24]) );
  dp_1 \pipeline/csr/mtvec_reg[25]  ( .ip(n9967), .ck(clk), .q(
        \pipeline/csr/mtvec [25]) );
  dp_1 \pipeline/csr/mtvec_reg[26]  ( .ip(n9966), .ck(clk), .q(
        \pipeline/csr/mtvec [26]) );
  dp_1 \pipeline/csr/mtvec_reg[27]  ( .ip(n9965), .ck(clk), .q(
        \pipeline/csr/mtvec [27]) );
  dp_1 \pipeline/csr/mtvec_reg[28]  ( .ip(n9964), .ck(clk), .q(
        \pipeline/csr/mtvec [28]) );
  dp_1 \pipeline/csr/mtvec_reg[29]  ( .ip(n9963), .ck(clk), .q(
        \pipeline/csr/mtvec [29]) );
  dp_1 \pipeline/csr/mtvec_reg[30]  ( .ip(n9962), .ck(clk), .q(
        \pipeline/csr/mtvec [30]) );
  dp_1 \pipeline/csr/mtvec_reg[31]  ( .ip(n9961), .ck(clk), .q(
        \pipeline/csr/mtvec [31]) );
  dp_1 \pipeline/csr/from_host_reg[0]  ( .ip(n9960), .ck(clk), .q(
        \pipeline/csr/from_host [0]) );
  dp_1 \pipeline/csr/from_host_reg[1]  ( .ip(n9959), .ck(clk), .q(
        \pipeline/csr/from_host [1]) );
  dp_1 \pipeline/csr/from_host_reg[2]  ( .ip(n9958), .ck(clk), .q(
        \pipeline/csr/from_host [2]) );
  dp_1 \pipeline/csr/from_host_reg[3]  ( .ip(n9957), .ck(clk), .q(
        \pipeline/csr/from_host [3]) );
  dp_1 \pipeline/csr/from_host_reg[4]  ( .ip(n9956), .ck(clk), .q(
        \pipeline/csr/from_host [4]) );
  dp_1 \pipeline/csr/from_host_reg[5]  ( .ip(n9955), .ck(clk), .q(
        \pipeline/csr/from_host [5]) );
  dp_1 \pipeline/csr/from_host_reg[6]  ( .ip(n9954), .ck(clk), .q(
        \pipeline/csr/from_host [6]) );
  dp_1 \pipeline/csr/from_host_reg[7]  ( .ip(n9953), .ck(clk), .q(
        \pipeline/csr/from_host [7]) );
  dp_1 \pipeline/csr/from_host_reg[8]  ( .ip(n9952), .ck(clk), .q(
        \pipeline/csr/from_host [8]) );
  dp_1 \pipeline/csr/from_host_reg[9]  ( .ip(n9951), .ck(clk), .q(
        \pipeline/csr/from_host [9]) );
  dp_1 \pipeline/csr/from_host_reg[10]  ( .ip(n9950), .ck(clk), .q(
        \pipeline/csr/from_host [10]) );
  dp_1 \pipeline/csr/from_host_reg[11]  ( .ip(n9949), .ck(clk), .q(
        \pipeline/csr/from_host [11]) );
  dp_1 \pipeline/csr/from_host_reg[12]  ( .ip(n9948), .ck(clk), .q(
        \pipeline/csr/from_host [12]) );
  dp_1 \pipeline/csr/from_host_reg[13]  ( .ip(n9947), .ck(clk), .q(
        \pipeline/csr/from_host [13]) );
  dp_1 \pipeline/csr/from_host_reg[14]  ( .ip(n9946), .ck(clk), .q(
        \pipeline/csr/from_host [14]) );
  dp_1 \pipeline/csr/from_host_reg[15]  ( .ip(n9945), .ck(clk), .q(
        \pipeline/csr/from_host [15]) );
  dp_1 \pipeline/csr/from_host_reg[16]  ( .ip(n9944), .ck(clk), .q(
        \pipeline/csr/from_host [16]) );
  dp_1 \pipeline/csr/from_host_reg[17]  ( .ip(n9943), .ck(clk), .q(
        \pipeline/csr/from_host [17]) );
  dp_1 \pipeline/csr/from_host_reg[18]  ( .ip(n9942), .ck(clk), .q(
        \pipeline/csr/from_host [18]) );
  dp_1 \pipeline/csr/from_host_reg[19]  ( .ip(n9941), .ck(clk), .q(
        \pipeline/csr/from_host [19]) );
  dp_1 \pipeline/csr/from_host_reg[20]  ( .ip(n9940), .ck(clk), .q(
        \pipeline/csr/from_host [20]) );
  dp_1 \pipeline/csr/from_host_reg[21]  ( .ip(n9939), .ck(clk), .q(
        \pipeline/csr/from_host [21]) );
  dp_1 \pipeline/csr/from_host_reg[22]  ( .ip(n9938), .ck(clk), .q(
        \pipeline/csr/from_host [22]) );
  dp_1 \pipeline/csr/from_host_reg[23]  ( .ip(n9937), .ck(clk), .q(
        \pipeline/csr/from_host [23]) );
  dp_1 \pipeline/csr/from_host_reg[24]  ( .ip(n9936), .ck(clk), .q(
        \pipeline/csr/from_host [24]) );
  dp_1 \pipeline/csr/from_host_reg[25]  ( .ip(n9935), .ck(clk), .q(
        \pipeline/csr/from_host [25]) );
  dp_1 \pipeline/csr/from_host_reg[26]  ( .ip(n9934), .ck(clk), .q(
        \pipeline/csr/from_host [26]) );
  dp_1 \pipeline/csr/from_host_reg[27]  ( .ip(n9933), .ck(clk), .q(
        \pipeline/csr/from_host [27]) );
  dp_1 \pipeline/csr/from_host_reg[28]  ( .ip(n9932), .ck(clk), .q(
        \pipeline/csr/from_host [28]) );
  dp_1 \pipeline/csr/from_host_reg[29]  ( .ip(n9931), .ck(clk), .q(
        \pipeline/csr/from_host [29]) );
  dp_1 \pipeline/csr/from_host_reg[30]  ( .ip(n9930), .ck(clk), .q(
        \pipeline/csr/from_host [30]) );
  dp_1 \pipeline/csr/from_host_reg[31]  ( .ip(n9929), .ck(clk), .q(
        \pipeline/csr/from_host [31]) );
  dp_1 \pipeline/csr/mscratch_reg[0]  ( .ip(n9928), .ck(clk), .q(
        \pipeline/csr/mscratch [0]) );
  dp_1 \pipeline/csr/mscratch_reg[1]  ( .ip(n9927), .ck(clk), .q(
        \pipeline/csr/mscratch [1]) );
  dp_1 \pipeline/csr/mscratch_reg[2]  ( .ip(n9926), .ck(clk), .q(
        \pipeline/csr/mscratch [2]) );
  dp_1 \pipeline/csr/mscratch_reg[3]  ( .ip(n9925), .ck(clk), .q(
        \pipeline/csr/mscratch [3]) );
  dp_1 \pipeline/csr/mscratch_reg[4]  ( .ip(n9924), .ck(clk), .q(
        \pipeline/csr/mscratch [4]) );
  dp_1 \pipeline/csr/mscratch_reg[5]  ( .ip(n9923), .ck(clk), .q(
        \pipeline/csr/mscratch [5]) );
  dp_1 \pipeline/csr/mscratch_reg[6]  ( .ip(n9922), .ck(clk), .q(
        \pipeline/csr/mscratch [6]) );
  dp_1 \pipeline/csr/mscratch_reg[7]  ( .ip(n9921), .ck(clk), .q(
        \pipeline/csr/mscratch [7]) );
  dp_1 \pipeline/csr/mscratch_reg[8]  ( .ip(n9920), .ck(clk), .q(
        \pipeline/csr/mscratch [8]) );
  dp_1 \pipeline/csr/mscratch_reg[9]  ( .ip(n9919), .ck(clk), .q(
        \pipeline/csr/mscratch [9]) );
  dp_1 \pipeline/csr/mscratch_reg[10]  ( .ip(n9918), .ck(clk), .q(
        \pipeline/csr/mscratch [10]) );
  dp_1 \pipeline/csr/mscratch_reg[11]  ( .ip(n9917), .ck(clk), .q(
        \pipeline/csr/mscratch [11]) );
  dp_1 \pipeline/csr/mscratch_reg[12]  ( .ip(n9916), .ck(clk), .q(
        \pipeline/csr/mscratch [12]) );
  dp_1 \pipeline/csr/mscratch_reg[13]  ( .ip(n9915), .ck(clk), .q(
        \pipeline/csr/mscratch [13]) );
  dp_1 \pipeline/csr/mscratch_reg[14]  ( .ip(n9914), .ck(clk), .q(
        \pipeline/csr/mscratch [14]) );
  dp_1 \pipeline/csr/mscratch_reg[15]  ( .ip(n9913), .ck(clk), .q(
        \pipeline/csr/mscratch [15]) );
  dp_1 \pipeline/csr/mscratch_reg[16]  ( .ip(n9912), .ck(clk), .q(
        \pipeline/csr/mscratch [16]) );
  dp_1 \pipeline/csr/mscratch_reg[17]  ( .ip(n9911), .ck(clk), .q(
        \pipeline/csr/mscratch [17]) );
  dp_1 \pipeline/csr/mscratch_reg[18]  ( .ip(n9910), .ck(clk), .q(
        \pipeline/csr/mscratch [18]) );
  dp_1 \pipeline/csr/mscratch_reg[19]  ( .ip(n9909), .ck(clk), .q(
        \pipeline/csr/mscratch [19]) );
  dp_1 \pipeline/csr/mscratch_reg[20]  ( .ip(n9908), .ck(clk), .q(
        \pipeline/csr/mscratch [20]) );
  dp_1 \pipeline/csr/mscratch_reg[21]  ( .ip(n9907), .ck(clk), .q(
        \pipeline/csr/mscratch [21]) );
  dp_1 \pipeline/csr/mscratch_reg[22]  ( .ip(n9906), .ck(clk), .q(
        \pipeline/csr/mscratch [22]) );
  dp_1 \pipeline/csr/mscratch_reg[23]  ( .ip(n9905), .ck(clk), .q(
        \pipeline/csr/mscratch [23]) );
  dp_1 \pipeline/csr/mscratch_reg[24]  ( .ip(n9904), .ck(clk), .q(
        \pipeline/csr/mscratch [24]) );
  dp_1 \pipeline/csr/mscratch_reg[25]  ( .ip(n9903), .ck(clk), .q(
        \pipeline/csr/mscratch [25]) );
  dp_1 \pipeline/csr/mscratch_reg[26]  ( .ip(n9902), .ck(clk), .q(
        \pipeline/csr/mscratch [26]) );
  dp_1 \pipeline/csr/mscratch_reg[27]  ( .ip(n9901), .ck(clk), .q(
        \pipeline/csr/mscratch [27]) );
  dp_1 \pipeline/csr/mscratch_reg[28]  ( .ip(n9900), .ck(clk), .q(
        \pipeline/csr/mscratch [28]) );
  dp_1 \pipeline/csr/mscratch_reg[29]  ( .ip(n9899), .ck(clk), .q(
        \pipeline/csr/mscratch [29]) );
  dp_1 \pipeline/csr/mscratch_reg[30]  ( .ip(n9898), .ck(clk), .q(
        \pipeline/csr/mscratch [30]) );
  dp_1 \pipeline/csr/mscratch_reg[31]  ( .ip(n9897), .ck(clk), .q(
        \pipeline/csr/mscratch [31]) );
  dp_1 \pipeline/csr/priv_stack_reg[5]  ( .ip(n10028), .ck(clk), .q(
        \pipeline/csr/priv_stack [5]) );
  dp_1 \pipeline/csr/priv_stack_reg[0]  ( .ip(n10027), .ck(clk), .q(
        \pipeline/csr/priv_stack_0 ) );
  dp_1 \pipeline/csr/priv_stack_reg[3]  ( .ip(n10024), .ck(clk), .q(
        \pipeline/csr/priv_stack [3]) );
  dp_1 \pipeline/csr/priv_stack_reg[4]  ( .ip(n10023), .ck(clk), .q(
        \pipeline/csr/priv_stack [4]) );
  dp_1 \pipeline/csr/mepc_reg[2]  ( .ip(n8869), .ck(clk), .q(\pipeline/epc [2]) );
  dp_1 \pipeline/csr/mepc_reg[3]  ( .ip(n8868), .ck(clk), .q(\pipeline/epc [3]) );
  dp_1 \pipeline/csr/mepc_reg[4]  ( .ip(n8867), .ck(clk), .q(\pipeline/epc [4]) );
  dp_1 \pipeline/csr/mepc_reg[5]  ( .ip(n8866), .ck(clk), .q(\pipeline/epc [5]) );
  dp_1 \pipeline/csr/mepc_reg[6]  ( .ip(n8865), .ck(clk), .q(\pipeline/epc [6]) );
  dp_1 \pipeline/csr/mepc_reg[7]  ( .ip(n8864), .ck(clk), .q(\pipeline/epc [7]) );
  dp_1 \pipeline/csr/mepc_reg[8]  ( .ip(n22851), .ck(clk), .q(
        \pipeline/epc [8]) );
  dp_1 \pipeline/csr/mepc_reg[9]  ( .ip(n8862), .ck(clk), .q(\pipeline/epc [9]) );
  dp_1 \pipeline/csr/mepc_reg[10]  ( .ip(n8861), .ck(clk), .q(
        \pipeline/epc [10]) );
  dp_1 \pipeline/csr/mepc_reg[11]  ( .ip(n22852), .ck(clk), .q(
        \pipeline/epc [11]) );
  dp_1 \pipeline/csr/mepc_reg[12]  ( .ip(n8859), .ck(clk), .q(
        \pipeline/epc [12]) );
  dp_1 \pipeline/csr/mepc_reg[13]  ( .ip(n8858), .ck(clk), .q(
        \pipeline/epc [13]) );
  dp_1 \pipeline/csr/mepc_reg[14]  ( .ip(n8857), .ck(clk), .q(
        \pipeline/epc [14]) );
  dp_1 \pipeline/csr/mepc_reg[15]  ( .ip(n8856), .ck(clk), .q(
        \pipeline/epc [15]) );
  dp_1 \pipeline/csr/mepc_reg[16]  ( .ip(n8855), .ck(clk), .q(
        \pipeline/epc [16]) );
  dp_1 \pipeline/csr/mepc_reg[17]  ( .ip(n8854), .ck(clk), .q(
        \pipeline/epc [17]) );
  dp_1 \pipeline/csr/mepc_reg[18]  ( .ip(n8853), .ck(clk), .q(
        \pipeline/epc [18]) );
  dp_1 \pipeline/csr/mepc_reg[19]  ( .ip(n8852), .ck(clk), .q(
        \pipeline/epc [19]) );
  dp_1 \pipeline/csr/mepc_reg[20]  ( .ip(n8851), .ck(clk), .q(
        \pipeline/epc [20]) );
  dp_1 \pipeline/csr/mepc_reg[21]  ( .ip(n8850), .ck(clk), .q(
        \pipeline/epc [21]) );
  dp_1 \pipeline/csr/mepc_reg[22]  ( .ip(n8849), .ck(clk), .q(
        \pipeline/epc [22]) );
  dp_1 \pipeline/csr/mepc_reg[23]  ( .ip(n8848), .ck(clk), .q(
        \pipeline/epc [23]) );
  dp_1 \pipeline/csr/mepc_reg[24]  ( .ip(n8847), .ck(clk), .q(
        \pipeline/epc [24]) );
  dp_1 \pipeline/csr/mepc_reg[25]  ( .ip(n8846), .ck(clk), .q(
        \pipeline/epc [25]) );
  dp_1 \pipeline/csr/mepc_reg[26]  ( .ip(n8845), .ck(clk), .q(
        \pipeline/epc [26]) );
  dp_1 \pipeline/csr/mepc_reg[27]  ( .ip(n8844), .ck(clk), .q(
        \pipeline/epc [27]) );
  dp_1 \pipeline/csr/mepc_reg[28]  ( .ip(n22863), .ck(clk), .q(
        \pipeline/epc [28]) );
  dp_1 \pipeline/csr/mepc_reg[29]  ( .ip(n8842), .ck(clk), .q(
        \pipeline/epc [29]) );
  dp_1 \pipeline/csr/mepc_reg[30]  ( .ip(n8841), .ck(clk), .q(
        \pipeline/epc [30]) );
  dp_1 \pipeline/csr/mepc_reg[31]  ( .ip(n8840), .ck(clk), .q(
        \pipeline/epc [31]) );
  dp_1 \pipeline/md/out_sel_reg[1]  ( .ip(n10063), .ck(clk), .q(
        \pipeline/md/out_sel [1]) );
  dp_1 \pipeline/md/out_sel_reg[0]  ( .ip(n10064), .ck(clk), .q(
        \pipeline/md/out_sel [0]) );
  dp_1 \pipeline/md/op_reg[0]  ( .ip(n10062), .ck(clk), .q(\pipeline/md/op [0]) );
  dp_1 \pipeline/md/op_reg[1]  ( .ip(n10061), .ck(clk), .q(\pipeline/md/op [1]) );
  dp_1 \pipeline/md/negate_output_reg  ( .ip(n8904), .ck(clk), .q(
        \pipeline/md/negate_output ) );
  dp_1 \pipeline/ctrl/prev_ex_code_WB_reg[3]  ( .ip(n8739), .ck(clk), .q(
        \pipeline/ctrl/prev_ex_code_WB [3]) );
  dp_1 \pipeline/ctrl/prev_ex_code_WB_reg[0]  ( .ip(n8738), .ck(clk), .q(
        \pipeline/ctrl/prev_ex_code_WB [0]) );
  dp_1 \pipeline/ctrl/prev_ex_code_WB_reg[1]  ( .ip(n8737), .ck(clk), .q(
        \pipeline/ctrl/prev_ex_code_WB [1]) );
  dp_1 \pipeline/csr/instret_full_reg[0]  ( .ip(n10138), .ck(clk), .q(
        \pipeline/csr/instret_full [0]) );
  dp_1 \pipeline/csr/instret_full_reg[1]  ( .ip(n10137), .ck(clk), .q(
        \pipeline/csr/instret_full [1]) );
  dp_1 \pipeline/csr/instret_full_reg[2]  ( .ip(n10136), .ck(clk), .q(
        \pipeline/csr/instret_full [2]) );
  dp_1 \pipeline/csr/instret_full_reg[3]  ( .ip(n10135), .ck(clk), .q(
        \pipeline/csr/instret_full [3]) );
  dp_1 \pipeline/csr/instret_full_reg[4]  ( .ip(n10134), .ck(clk), .q(
        \pipeline/csr/instret_full [4]) );
  dp_1 \pipeline/csr/instret_full_reg[5]  ( .ip(n10133), .ck(clk), .q(
        \pipeline/csr/instret_full [5]) );
  dp_1 \pipeline/csr/instret_full_reg[6]  ( .ip(n10132), .ck(clk), .q(
        \pipeline/csr/instret_full [6]) );
  dp_1 \pipeline/csr/instret_full_reg[7]  ( .ip(n10131), .ck(clk), .q(
        \pipeline/csr/instret_full [7]) );
  dp_1 \pipeline/csr/instret_full_reg[8]  ( .ip(n22858), .ck(clk), .q(
        \pipeline/csr/instret_full [8]) );
  dp_1 \pipeline/csr/instret_full_reg[9]  ( .ip(n10129), .ck(clk), .q(
        \pipeline/csr/instret_full [9]) );
  dp_1 \pipeline/csr/instret_full_reg[10]  ( .ip(n10128), .ck(clk), .q(
        \pipeline/csr/instret_full [10]) );
  dp_1 \pipeline/csr/instret_full_reg[11]  ( .ip(n22856), .ck(clk), .q(
        \pipeline/csr/instret_full [11]) );
  dp_1 \pipeline/csr/instret_full_reg[12]  ( .ip(n10126), .ck(clk), .q(
        \pipeline/csr/instret_full [12]) );
  dp_1 \pipeline/csr/instret_full_reg[13]  ( .ip(n10125), .ck(clk), .q(
        \pipeline/csr/instret_full [13]) );
  dp_1 \pipeline/csr/instret_full_reg[14]  ( .ip(n10124), .ck(clk), .q(
        \pipeline/csr/instret_full [14]) );
  dp_1 \pipeline/csr/instret_full_reg[15]  ( .ip(n10123), .ck(clk), .q(
        \pipeline/csr/instret_full [15]) );
  dp_1 \pipeline/csr/instret_full_reg[16]  ( .ip(n10122), .ck(clk), .q(
        \pipeline/csr/instret_full [16]) );
  dp_1 \pipeline/csr/instret_full_reg[17]  ( .ip(n10121), .ck(clk), .q(
        \pipeline/csr/instret_full [17]) );
  dp_1 \pipeline/csr/instret_full_reg[18]  ( .ip(n10120), .ck(clk), .q(
        \pipeline/csr/instret_full [18]) );
  dp_1 \pipeline/csr/instret_full_reg[19]  ( .ip(n10119), .ck(clk), .q(
        \pipeline/csr/instret_full [19]) );
  dp_1 \pipeline/csr/instret_full_reg[20]  ( .ip(n10118), .ck(clk), .q(
        \pipeline/csr/instret_full [20]) );
  dp_1 \pipeline/csr/instret_full_reg[21]  ( .ip(n10117), .ck(clk), .q(
        \pipeline/csr/instret_full [21]) );
  dp_1 \pipeline/csr/instret_full_reg[22]  ( .ip(n10116), .ck(clk), .q(
        \pipeline/csr/instret_full [22]) );
  dp_1 \pipeline/csr/instret_full_reg[23]  ( .ip(n10115), .ck(clk), .q(
        \pipeline/csr/instret_full [23]) );
  dp_1 \pipeline/csr/instret_full_reg[24]  ( .ip(n10114), .ck(clk), .q(
        \pipeline/csr/instret_full [24]) );
  dp_1 \pipeline/csr/instret_full_reg[25]  ( .ip(n10113), .ck(clk), .q(
        \pipeline/csr/instret_full [25]) );
  dp_1 \pipeline/csr/instret_full_reg[26]  ( .ip(n10112), .ck(clk), .q(
        \pipeline/csr/instret_full [26]) );
  dp_1 \pipeline/csr/instret_full_reg[27]  ( .ip(n10111), .ck(clk), .q(
        \pipeline/csr/instret_full [27]) );
  dp_1 \pipeline/csr/instret_full_reg[28]  ( .ip(n10110), .ck(clk), .q(
        \pipeline/csr/instret_full [28]) );
  dp_1 \pipeline/csr/instret_full_reg[29]  ( .ip(n10109), .ck(clk), .q(
        \pipeline/csr/instret_full [29]) );
  dp_1 \pipeline/csr/instret_full_reg[30]  ( .ip(n10108), .ck(clk), .q(
        \pipeline/csr/instret_full [30]) );
  dp_1 \pipeline/csr/instret_full_reg[31]  ( .ip(n10107), .ck(clk), .q(
        \pipeline/csr/instret_full [31]) );
  dp_1 \pipeline/csr/instret_full_reg[32]  ( .ip(n10106), .ck(clk), .q(
        \pipeline/csr/instret_full [32]) );
  dp_1 \pipeline/csr/instret_full_reg[33]  ( .ip(n10105), .ck(clk), .q(
        \pipeline/csr/instret_full [33]) );
  dp_1 \pipeline/csr/instret_full_reg[34]  ( .ip(n10104), .ck(clk), .q(
        \pipeline/csr/instret_full [34]) );
  dp_1 \pipeline/csr/instret_full_reg[35]  ( .ip(n10103), .ck(clk), .q(
        \pipeline/csr/instret_full [35]) );
  dp_1 \pipeline/csr/instret_full_reg[36]  ( .ip(n10102), .ck(clk), .q(
        \pipeline/csr/instret_full [36]) );
  dp_1 \pipeline/csr/instret_full_reg[37]  ( .ip(n10101), .ck(clk), .q(
        \pipeline/csr/instret_full [37]) );
  dp_1 \pipeline/csr/instret_full_reg[38]  ( .ip(n10100), .ck(clk), .q(
        \pipeline/csr/instret_full [38]) );
  dp_1 \pipeline/csr/instret_full_reg[39]  ( .ip(n10099), .ck(clk), .q(
        \pipeline/csr/instret_full [39]) );
  dp_1 \pipeline/csr/instret_full_reg[40]  ( .ip(n10098), .ck(clk), .q(
        \pipeline/csr/instret_full [40]) );
  dp_1 \pipeline/csr/instret_full_reg[41]  ( .ip(n10097), .ck(clk), .q(
        \pipeline/csr/instret_full [41]) );
  dp_1 \pipeline/csr/instret_full_reg[42]  ( .ip(n10096), .ck(clk), .q(
        \pipeline/csr/instret_full [42]) );
  dp_1 \pipeline/csr/instret_full_reg[43]  ( .ip(n22853), .ck(clk), .q(
        \pipeline/csr/instret_full [43]) );
  dp_1 \pipeline/csr/instret_full_reg[44]  ( .ip(n10094), .ck(clk), .q(
        \pipeline/csr/instret_full [44]) );
  dp_1 \pipeline/csr/instret_full_reg[45]  ( .ip(n10093), .ck(clk), .q(
        \pipeline/csr/instret_full [45]) );
  dp_1 \pipeline/csr/instret_full_reg[46]  ( .ip(n10092), .ck(clk), .q(
        \pipeline/csr/instret_full [46]) );
  dp_1 \pipeline/csr/instret_full_reg[47]  ( .ip(n10091), .ck(clk), .q(
        \pipeline/csr/instret_full [47]) );
  dp_1 \pipeline/csr/instret_full_reg[48]  ( .ip(n10090), .ck(clk), .q(
        \pipeline/csr/instret_full [48]) );
  dp_1 \pipeline/csr/instret_full_reg[49]  ( .ip(n10089), .ck(clk), .q(
        \pipeline/csr/instret_full [49]) );
  dp_1 \pipeline/csr/instret_full_reg[50]  ( .ip(n10088), .ck(clk), .q(
        \pipeline/csr/instret_full [50]) );
  dp_1 \pipeline/csr/instret_full_reg[51]  ( .ip(n10087), .ck(clk), .q(
        \pipeline/csr/instret_full [51]) );
  dp_1 \pipeline/csr/instret_full_reg[52]  ( .ip(n10086), .ck(clk), .q(
        \pipeline/csr/instret_full [52]) );
  dp_1 \pipeline/csr/instret_full_reg[53]  ( .ip(n10085), .ck(clk), .q(
        \pipeline/csr/instret_full [53]) );
  dp_1 \pipeline/csr/instret_full_reg[54]  ( .ip(n10084), .ck(clk), .q(
        \pipeline/csr/instret_full [54]) );
  dp_1 \pipeline/csr/instret_full_reg[55]  ( .ip(n10083), .ck(clk), .q(
        \pipeline/csr/instret_full [55]) );
  dp_1 \pipeline/csr/instret_full_reg[56]  ( .ip(n10082), .ck(clk), .q(
        \pipeline/csr/instret_full [56]) );
  dp_1 \pipeline/csr/instret_full_reg[57]  ( .ip(n10081), .ck(clk), .q(
        \pipeline/csr/instret_full [57]) );
  dp_1 \pipeline/csr/instret_full_reg[58]  ( .ip(n10080), .ck(clk), .q(
        \pipeline/csr/instret_full [58]) );
  dp_1 \pipeline/csr/instret_full_reg[59]  ( .ip(n10079), .ck(clk), .q(
        \pipeline/csr/instret_full [59]) );
  dp_1 \pipeline/csr/instret_full_reg[60]  ( .ip(n10078), .ck(clk), .q(
        \pipeline/csr/instret_full [60]) );
  dp_1 \pipeline/csr/instret_full_reg[61]  ( .ip(n10077), .ck(clk), .q(
        \pipeline/csr/instret_full [61]) );
  dp_1 \pipeline/csr/instret_full_reg[62]  ( .ip(n10076), .ck(clk), .q(
        \pipeline/csr/instret_full [62]) );
  dp_1 \pipeline/csr/instret_full_reg[63]  ( .ip(n10075), .ck(clk), .q(
        \pipeline/csr/instret_full [63]) );
  dp_1 \pipeline/csr/mint_reg  ( .ip(n8736), .ck(clk), .q(
        \pipeline/csr/mcause[31] ) );
  dp_1 \pipeline/csr/mecode_reg[0]  ( .ip(n8735), .ck(clk), .q(
        \pipeline/csr/mecode [0]) );
  dp_1 \pipeline/csr/mecode_reg[1]  ( .ip(n8734), .ck(clk), .q(
        \pipeline/csr/mecode [1]) );
  dp_1 \pipeline/csr/mecode_reg[2]  ( .ip(n8733), .ck(clk), .q(
        \pipeline/csr/mecode [2]) );
  dp_1 \pipeline/csr/mecode_reg[3]  ( .ip(n8732), .ck(clk), .q(
        \pipeline/csr/mecode [3]) );
  dp_1 \pipeline/PC_WB_reg[0]  ( .ip(n8903), .ck(clk), .q(\pipeline/PC_WB [0])
         );
  dp_1 \pipeline/PC_WB_reg[1]  ( .ip(n8902), .ck(clk), .q(\pipeline/PC_WB [1])
         );
  dp_1 \pipeline/PC_WB_reg[2]  ( .ip(n8901), .ck(clk), .q(\pipeline/PC_WB [2])
         );
  dp_1 \pipeline/PC_WB_reg[3]  ( .ip(n8900), .ck(clk), .q(\pipeline/PC_WB [3])
         );
  dp_1 \pipeline/PC_WB_reg[4]  ( .ip(n8899), .ck(clk), .q(\pipeline/PC_WB [4])
         );
  dp_1 \pipeline/PC_WB_reg[5]  ( .ip(n8898), .ck(clk), .q(\pipeline/PC_WB [5])
         );
  dp_1 \pipeline/PC_WB_reg[6]  ( .ip(n8897), .ck(clk), .q(\pipeline/PC_WB [6])
         );
  dp_1 \pipeline/PC_WB_reg[7]  ( .ip(n8896), .ck(clk), .q(\pipeline/PC_WB [7])
         );
  dp_1 \pipeline/PC_WB_reg[8]  ( .ip(n8895), .ck(clk), .q(\pipeline/PC_WB [8])
         );
  dp_1 \pipeline/PC_WB_reg[9]  ( .ip(n8894), .ck(clk), .q(\pipeline/PC_WB [9])
         );
  dp_1 \pipeline/PC_WB_reg[10]  ( .ip(n8893), .ck(clk), .q(
        \pipeline/PC_WB [10]) );
  dp_1 \pipeline/PC_WB_reg[11]  ( .ip(n8892), .ck(clk), .q(
        \pipeline/PC_WB [11]) );
  dp_1 \pipeline/PC_WB_reg[12]  ( .ip(n8891), .ck(clk), .q(
        \pipeline/PC_WB [12]) );
  dp_1 \pipeline/PC_WB_reg[13]  ( .ip(n8890), .ck(clk), .q(
        \pipeline/PC_WB [13]) );
  dp_1 \pipeline/PC_WB_reg[14]  ( .ip(n8889), .ck(clk), .q(
        \pipeline/PC_WB [14]) );
  dp_1 \pipeline/PC_WB_reg[15]  ( .ip(n8888), .ck(clk), .q(
        \pipeline/PC_WB [15]) );
  dp_1 \pipeline/PC_WB_reg[16]  ( .ip(n8887), .ck(clk), .q(
        \pipeline/PC_WB [16]) );
  dp_1 \pipeline/PC_WB_reg[17]  ( .ip(n8886), .ck(clk), .q(
        \pipeline/PC_WB [17]) );
  dp_1 \pipeline/PC_WB_reg[18]  ( .ip(n8885), .ck(clk), .q(
        \pipeline/PC_WB [18]) );
  dp_1 \pipeline/PC_WB_reg[19]  ( .ip(n8884), .ck(clk), .q(
        \pipeline/PC_WB [19]) );
  dp_1 \pipeline/PC_WB_reg[20]  ( .ip(n8883), .ck(clk), .q(
        \pipeline/PC_WB [20]) );
  dp_1 \pipeline/PC_WB_reg[21]  ( .ip(n8882), .ck(clk), .q(
        \pipeline/PC_WB [21]) );
  dp_1 \pipeline/PC_WB_reg[22]  ( .ip(n8881), .ck(clk), .q(
        \pipeline/PC_WB [22]) );
  dp_1 \pipeline/PC_WB_reg[23]  ( .ip(n8880), .ck(clk), .q(
        \pipeline/PC_WB [23]) );
  dp_1 \pipeline/PC_WB_reg[24]  ( .ip(n8879), .ck(clk), .q(
        \pipeline/PC_WB [24]) );
  dp_1 \pipeline/PC_WB_reg[25]  ( .ip(n8878), .ck(clk), .q(
        \pipeline/PC_WB [25]) );
  dp_1 \pipeline/PC_WB_reg[26]  ( .ip(n8877), .ck(clk), .q(
        \pipeline/PC_WB [26]) );
  dp_1 \pipeline/PC_WB_reg[27]  ( .ip(n8876), .ck(clk), .q(
        \pipeline/PC_WB [27]) );
  dp_1 \pipeline/PC_WB_reg[28]  ( .ip(n8875), .ck(clk), .q(
        \pipeline/PC_WB [28]) );
  dp_1 \pipeline/PC_WB_reg[29]  ( .ip(n8874), .ck(clk), .q(
        \pipeline/PC_WB [29]) );
  dp_1 \pipeline/PC_WB_reg[30]  ( .ip(n8873), .ck(clk), .q(
        \pipeline/PC_WB [30]) );
  dp_1 \pipeline/PC_WB_reg[31]  ( .ip(n8872), .ck(clk), .q(
        \pipeline/PC_WB [31]) );
  dp_1 \pipeline/alu_out_WB_reg[0]  ( .ip(n8807), .ck(clk), .q(
        \pipeline/alu_out_WB [0]) );
  dp_1 \pipeline/csr/mbadaddr_reg[0]  ( .ip(n8700), .ck(clk), .q(
        \pipeline/csr/mbadaddr [0]) );
  dp_1 \pipeline/csr_rdata_WB_reg[0]  ( .ip(n8806), .ck(clk), .q(
        \pipeline/csr_rdata_WB [0]) );
  dp_1 \pipeline/alu_out_WB_reg[16]  ( .ip(n8716), .ck(clk), .q(
        \pipeline/alu_out_WB [16]) );
  dp_1 \pipeline/csr/mbadaddr_reg[16]  ( .ip(n8684), .ck(clk), .q(
        \pipeline/csr/mbadaddr [16]) );
  dp_1 \pipeline/csr_rdata_WB_reg[16]  ( .ip(n8790), .ck(clk), .q(
        \pipeline/csr_rdata_WB [16]) );
  dp_1 \pipeline/store_data_WB_reg[16]  ( .ip(n8823), .ck(clk), .q(
        \pipeline/store_data_WB [16]) );
  dp_1 \pipeline/alu_out_WB_reg[24]  ( .ip(n8708), .ck(clk), .q(
        \pipeline/alu_out_WB [24]) );
  dp_1 \pipeline/csr/mbadaddr_reg[24]  ( .ip(n8676), .ck(clk), .q(
        \pipeline/csr/mbadaddr [24]) );
  dp_1 \pipeline/csr_rdata_WB_reg[24]  ( .ip(n8782), .ck(clk), .q(
        \pipeline/csr_rdata_WB [24]) );
  dp_1 \pipeline/store_data_WB_reg[24]  ( .ip(n8815), .ck(clk), .q(
        \pipeline/store_data_WB [24]) );
  dp_1 \pipeline/alu_out_WB_reg[28]  ( .ip(n8704), .ck(clk), .q(
        \pipeline/alu_out_WB [28]) );
  dp_1 \pipeline/csr/mbadaddr_reg[28]  ( .ip(n8672), .ck(clk), .q(
        \pipeline/csr/mbadaddr [28]) );
  dp_1 \pipeline/csr_rdata_WB_reg[28]  ( .ip(n8778), .ck(clk), .q(
        \pipeline/csr_rdata_WB [28]) );
  dp_1 \pipeline/store_data_WB_reg[28]  ( .ip(n8811), .ck(clk), .q(
        \pipeline/store_data_WB [28]) );
  dp_1 \pipeline/alu_out_WB_reg[30]  ( .ip(n8702), .ck(clk), .q(
        \pipeline/alu_out_WB [30]) );
  dp_1 \pipeline/csr/mbadaddr_reg[30]  ( .ip(n8670), .ck(clk), .q(
        \pipeline/csr/mbadaddr [30]) );
  dp_1 \pipeline/csr_rdata_WB_reg[30]  ( .ip(n8776), .ck(clk), .q(
        \pipeline/csr_rdata_WB [30]) );
  dp_1 \pipeline/store_data_WB_reg[30]  ( .ip(n8809), .ck(clk), .q(
        \pipeline/store_data_WB [30]) );
  dp_1 \pipeline/alu_out_WB_reg[11]  ( .ip(n8721), .ck(clk), .q(
        \pipeline/alu_out_WB [11]) );
  dp_1 \pipeline/csr/mbadaddr_reg[11]  ( .ip(n8689), .ck(clk), .q(
        \pipeline/csr/mbadaddr [11]) );
  dp_1 \pipeline/csr_rdata_WB_reg[11]  ( .ip(n8795), .ck(clk), .q(
        \pipeline/csr_rdata_WB [11]) );
  dp_1 \pipeline/store_data_WB_reg[11]  ( .ip(n8828), .ck(clk), .q(
        \pipeline/store_data_WB [11]) );
  dp_1 \pipeline/alu_out_WB_reg[27]  ( .ip(n8705), .ck(clk), .q(
        \pipeline/alu_out_WB [27]) );
  dp_1 \pipeline/csr/mbadaddr_reg[27]  ( .ip(n8673), .ck(clk), .q(
        \pipeline/csr/mbadaddr [27]) );
  dp_1 \pipeline/csr_rdata_WB_reg[27]  ( .ip(n8779), .ck(clk), .q(
        \pipeline/csr_rdata_WB [27]) );
  dp_1 \pipeline/store_data_WB_reg[27]  ( .ip(n8812), .ck(clk), .q(
        \pipeline/store_data_WB [27]) );
  dp_1 \pipeline/alu_out_WB_reg[29]  ( .ip(n8703), .ck(clk), .q(
        \pipeline/alu_out_WB [29]) );
  dp_1 \pipeline/csr/mbadaddr_reg[29]  ( .ip(n8671), .ck(clk), .q(
        \pipeline/csr/mbadaddr [29]) );
  dp_1 \pipeline/csr_rdata_WB_reg[29]  ( .ip(n8777), .ck(clk), .q(
        \pipeline/csr_rdata_WB [29]) );
  dp_1 \pipeline/store_data_WB_reg[29]  ( .ip(n8810), .ck(clk), .q(
        \pipeline/store_data_WB [29]) );
  dp_1 \pipeline/alu_out_WB_reg[10]  ( .ip(n8722), .ck(clk), .q(
        \pipeline/alu_out_WB [10]) );
  dp_1 \pipeline/csr/mbadaddr_reg[10]  ( .ip(n8690), .ck(clk), .q(
        \pipeline/csr/mbadaddr [10]) );
  dp_1 \pipeline/csr_rdata_WB_reg[10]  ( .ip(n8796), .ck(clk), .q(
        \pipeline/csr_rdata_WB [10]) );
  dp_1 \pipeline/store_data_WB_reg[10]  ( .ip(n8829), .ck(clk), .q(
        \pipeline/store_data_WB [10]) );
  dp_1 \pipeline/alu_out_WB_reg[26]  ( .ip(n8706), .ck(clk), .q(
        \pipeline/alu_out_WB [26]) );
  dp_1 \pipeline/csr/mbadaddr_reg[26]  ( .ip(n8674), .ck(clk), .q(
        \pipeline/csr/mbadaddr [26]) );
  dp_1 \pipeline/csr_rdata_WB_reg[26]  ( .ip(n8780), .ck(clk), .q(
        \pipeline/csr_rdata_WB [26]) );
  dp_1 \pipeline/store_data_WB_reg[26]  ( .ip(n8813), .ck(clk), .q(
        \pipeline/store_data_WB [26]) );
  dp_1 \pipeline/alu_out_WB_reg[12]  ( .ip(n8720), .ck(clk), .q(
        \pipeline/alu_out_WB [12]) );
  dp_1 \pipeline/csr/mbadaddr_reg[12]  ( .ip(n8688), .ck(clk), .q(
        \pipeline/csr/mbadaddr [12]) );
  dp_1 \pipeline/csr_rdata_WB_reg[12]  ( .ip(n8794), .ck(clk), .q(
        \pipeline/csr_rdata_WB [12]) );
  dp_1 \pipeline/store_data_WB_reg[12]  ( .ip(n8827), .ck(clk), .q(
        \pipeline/store_data_WB [12]) );
  dp_1 \pipeline/alu_out_WB_reg[20]  ( .ip(n8712), .ck(clk), .q(
        \pipeline/alu_out_WB [20]) );
  dp_1 \pipeline/csr/mbadaddr_reg[20]  ( .ip(n8680), .ck(clk), .q(
        \pipeline/csr/mbadaddr [20]) );
  dp_1 \pipeline/csr_rdata_WB_reg[20]  ( .ip(n8786), .ck(clk), .q(
        \pipeline/csr_rdata_WB [20]) );
  dp_1 \pipeline/store_data_WB_reg[20]  ( .ip(n8819), .ck(clk), .q(
        \pipeline/store_data_WB [20]) );
  dp_1 \pipeline/alu_out_WB_reg[22]  ( .ip(n8710), .ck(clk), .q(
        \pipeline/alu_out_WB [22]) );
  dp_1 \pipeline/csr/mbadaddr_reg[22]  ( .ip(n8678), .ck(clk), .q(
        \pipeline/csr/mbadaddr [22]) );
  dp_1 \pipeline/csr_rdata_WB_reg[22]  ( .ip(n8784), .ck(clk), .q(
        \pipeline/csr_rdata_WB [22]) );
  dp_1 \pipeline/store_data_WB_reg[22]  ( .ip(n8817), .ck(clk), .q(
        \pipeline/store_data_WB [22]) );
  dp_1 \pipeline/alu_out_WB_reg[23]  ( .ip(n8709), .ck(clk), .q(
        \pipeline/alu_out_WB [23]) );
  dp_1 \pipeline/csr/mbadaddr_reg[23]  ( .ip(n8677), .ck(clk), .q(
        \pipeline/csr/mbadaddr [23]) );
  dp_1 \pipeline/csr_rdata_WB_reg[23]  ( .ip(n8783), .ck(clk), .q(
        \pipeline/csr_rdata_WB [23]) );
  dp_1 \pipeline/store_data_WB_reg[23]  ( .ip(n8816), .ck(clk), .q(
        \pipeline/store_data_WB [23]) );
  dp_1 \pipeline/alu_out_WB_reg[8]  ( .ip(n8724), .ck(clk), .q(
        \pipeline/alu_out_WB [8]) );
  dp_1 \pipeline/csr/mbadaddr_reg[8]  ( .ip(n8692), .ck(clk), .q(
        \pipeline/csr/mbadaddr [8]) );
  dp_1 \pipeline/csr_rdata_WB_reg[8]  ( .ip(n8798), .ck(clk), .q(
        \pipeline/csr_rdata_WB [8]) );
  dp_1 \pipeline/store_data_WB_reg[8]  ( .ip(n8831), .ck(clk), .q(
        \pipeline/store_data_WB [8]) );
  dp_1 \pipeline/alu_out_WB_reg[13]  ( .ip(n8719), .ck(clk), .q(
        \pipeline/alu_out_WB [13]) );
  dp_1 \pipeline/csr/mbadaddr_reg[13]  ( .ip(n8687), .ck(clk), .q(
        \pipeline/csr/mbadaddr [13]) );
  dp_1 \pipeline/csr_rdata_WB_reg[13]  ( .ip(n8793), .ck(clk), .q(
        \pipeline/csr_rdata_WB [13]) );
  dp_1 \pipeline/store_data_WB_reg[13]  ( .ip(n8826), .ck(clk), .q(
        \pipeline/store_data_WB [13]) );
  dp_1 \pipeline/alu_out_WB_reg[17]  ( .ip(n8715), .ck(clk), .q(
        \pipeline/alu_out_WB [17]) );
  dp_1 \pipeline/csr/mbadaddr_reg[17]  ( .ip(n8683), .ck(clk), .q(
        \pipeline/csr/mbadaddr [17]) );
  dp_1 \pipeline/csr_rdata_WB_reg[17]  ( .ip(n8789), .ck(clk), .q(
        \pipeline/csr_rdata_WB [17]) );
  dp_1 \pipeline/store_data_WB_reg[17]  ( .ip(n8822), .ck(clk), .q(
        \pipeline/store_data_WB [17]) );
  dp_1 \pipeline/alu_out_WB_reg[21]  ( .ip(n8711), .ck(clk), .q(
        \pipeline/alu_out_WB [21]) );
  dp_1 \pipeline/csr/mbadaddr_reg[21]  ( .ip(n8679), .ck(clk), .q(
        \pipeline/csr/mbadaddr [21]) );
  dp_1 \pipeline/csr_rdata_WB_reg[21]  ( .ip(n8785), .ck(clk), .q(
        \pipeline/csr_rdata_WB [21]) );
  dp_1 \pipeline/store_data_WB_reg[21]  ( .ip(n8818), .ck(clk), .q(
        \pipeline/store_data_WB [21]) );
  dp_1 \pipeline/alu_out_WB_reg[25]  ( .ip(n8707), .ck(clk), .q(
        \pipeline/alu_out_WB [25]) );
  dp_1 \pipeline/csr/mbadaddr_reg[25]  ( .ip(n8675), .ck(clk), .q(
        \pipeline/csr/mbadaddr [25]) );
  dp_1 \pipeline/csr_rdata_WB_reg[25]  ( .ip(n8781), .ck(clk), .q(
        \pipeline/csr_rdata_WB [25]) );
  dp_1 \pipeline/store_data_WB_reg[25]  ( .ip(n8814), .ck(clk), .q(
        \pipeline/store_data_WB [25]) );
  dp_1 \pipeline/alu_out_WB_reg[18]  ( .ip(n8714), .ck(clk), .q(
        \pipeline/alu_out_WB [18]) );
  dp_1 \pipeline/csr/mbadaddr_reg[18]  ( .ip(n8682), .ck(clk), .q(
        \pipeline/csr/mbadaddr [18]) );
  dp_1 \pipeline/csr_rdata_WB_reg[18]  ( .ip(n8788), .ck(clk), .q(
        \pipeline/csr_rdata_WB [18]) );
  dp_1 \pipeline/store_data_WB_reg[18]  ( .ip(n8821), .ck(clk), .q(
        \pipeline/store_data_WB [18]) );
  dp_1 \pipeline/alu_out_WB_reg[19]  ( .ip(n8713), .ck(clk), .q(
        \pipeline/alu_out_WB [19]) );
  dp_1 \pipeline/csr/mbadaddr_reg[19]  ( .ip(n8681), .ck(clk), .q(
        \pipeline/csr/mbadaddr [19]) );
  dp_1 \pipeline/csr_rdata_WB_reg[19]  ( .ip(n8787), .ck(clk), .q(
        \pipeline/csr_rdata_WB [19]) );
  dp_1 \pipeline/store_data_WB_reg[19]  ( .ip(n8820), .ck(clk), .q(
        \pipeline/store_data_WB [19]) );
  dp_1 \pipeline/alu_out_WB_reg[4]  ( .ip(n8728), .ck(clk), .q(
        \pipeline/alu_out_WB [4]) );
  dp_1 \pipeline/csr/mbadaddr_reg[4]  ( .ip(n8696), .ck(clk), .q(
        \pipeline/csr/mbadaddr [4]) );
  dp_1 \pipeline/csr_rdata_WB_reg[4]  ( .ip(n8802), .ck(clk), .q(
        \pipeline/csr_rdata_WB [4]) );
  dp_1 \pipeline/store_data_WB_reg[4]  ( .ip(n8835), .ck(clk), .q(
        dmem_hwdata[4]) );
  dp_1 \pipeline/alu_out_WB_reg[14]  ( .ip(n8718), .ck(clk), .q(
        \pipeline/alu_out_WB [14]) );
  dp_1 \pipeline/csr/mbadaddr_reg[14]  ( .ip(n8686), .ck(clk), .q(
        \pipeline/csr/mbadaddr [14]) );
  dp_1 \pipeline/csr_rdata_WB_reg[14]  ( .ip(n8792), .ck(clk), .q(
        \pipeline/csr_rdata_WB [14]) );
  dp_1 \pipeline/store_data_WB_reg[14]  ( .ip(n8825), .ck(clk), .q(
        \pipeline/store_data_WB [14]) );
  dp_1 \pipeline/alu_out_WB_reg[15]  ( .ip(n8717), .ck(clk), .q(
        \pipeline/alu_out_WB [15]) );
  dp_1 \pipeline/csr/mbadaddr_reg[15]  ( .ip(n8685), .ck(clk), .q(
        \pipeline/csr/mbadaddr [15]) );
  dp_1 \pipeline/csr_rdata_WB_reg[15]  ( .ip(n8791), .ck(clk), .q(
        \pipeline/csr_rdata_WB [15]) );
  dp_1 \pipeline/store_data_WB_reg[15]  ( .ip(n8824), .ck(clk), .q(
        \pipeline/store_data_WB [15]) );
  dp_1 \pipeline/alu_out_WB_reg[2]  ( .ip(n8730), .ck(clk), .q(
        \pipeline/alu_out_WB [2]) );
  dp_1 \pipeline/csr/mbadaddr_reg[2]  ( .ip(n8698), .ck(clk), .q(
        \pipeline/csr/mbadaddr [2]) );
  dp_1 \pipeline/csr_rdata_WB_reg[2]  ( .ip(n8804), .ck(clk), .q(
        \pipeline/csr_rdata_WB [2]) );
  dp_1 \pipeline/store_data_WB_reg[2]  ( .ip(n8837), .ck(clk), .q(
        dmem_hwdata[2]) );
  dp_1 \pipeline/alu_out_WB_reg[3]  ( .ip(n8729), .ck(clk), .q(
        \pipeline/alu_out_WB [3]) );
  dp_1 \pipeline/csr/mbadaddr_reg[3]  ( .ip(n8697), .ck(clk), .q(
        \pipeline/csr/mbadaddr [3]) );
  dp_1 \pipeline/csr_rdata_WB_reg[3]  ( .ip(n8803), .ck(clk), .q(
        \pipeline/csr_rdata_WB [3]) );
  dp_1 \pipeline/store_data_WB_reg[3]  ( .ip(n8836), .ck(clk), .q(
        dmem_hwdata[3]) );
  dp_1 \pipeline/alu_out_WB_reg[1]  ( .ip(n8731), .ck(clk), .q(
        \pipeline/alu_out_WB [1]) );
  dp_1 \pipeline/csr/mbadaddr_reg[1]  ( .ip(n8699), .ck(clk), .q(
        \pipeline/csr/mbadaddr [1]) );
  dp_1 \pipeline/csr_rdata_WB_reg[1]  ( .ip(n8805), .ck(clk), .q(
        \pipeline/csr_rdata_WB [1]) );
  dp_1 \pipeline/store_data_WB_reg[1]  ( .ip(n8838), .ck(clk), .q(
        dmem_hwdata[1]) );
  dp_1 \pipeline/alu_out_WB_reg[5]  ( .ip(n8727), .ck(clk), .q(
        \pipeline/alu_out_WB [5]) );
  dp_1 \pipeline/csr/mbadaddr_reg[5]  ( .ip(n8695), .ck(clk), .q(
        \pipeline/csr/mbadaddr [5]) );
  dp_1 \pipeline/csr_rdata_WB_reg[5]  ( .ip(n8801), .ck(clk), .q(
        \pipeline/csr_rdata_WB [5]) );
  dp_1 \pipeline/store_data_WB_reg[5]  ( .ip(n8834), .ck(clk), .q(
        dmem_hwdata[5]) );
  dp_1 \pipeline/alu_out_WB_reg[9]  ( .ip(n8723), .ck(clk), .q(
        \pipeline/alu_out_WB [9]) );
  dp_1 \pipeline/csr/mbadaddr_reg[9]  ( .ip(n8691), .ck(clk), .q(
        \pipeline/csr/mbadaddr [9]) );
  dp_1 \pipeline/csr_rdata_WB_reg[9]  ( .ip(n8797), .ck(clk), .q(
        \pipeline/csr_rdata_WB [9]) );
  dp_1 \pipeline/store_data_WB_reg[9]  ( .ip(n8830), .ck(clk), .q(
        \pipeline/store_data_WB [9]) );
  dp_1 \pipeline/alu_out_WB_reg[7]  ( .ip(n8725), .ck(clk), .q(
        \pipeline/alu_out_WB [7]) );
  dp_1 \pipeline/csr/mbadaddr_reg[7]  ( .ip(n8693), .ck(clk), .q(
        \pipeline/csr/mbadaddr [7]) );
  dp_1 \pipeline/csr_rdata_WB_reg[7]  ( .ip(n8799), .ck(clk), .q(
        \pipeline/csr_rdata_WB [7]) );
  dp_1 \pipeline/store_data_WB_reg[7]  ( .ip(n8832), .ck(clk), .q(
        dmem_hwdata[7]) );
  dp_1 \pipeline/alu_out_WB_reg[6]  ( .ip(n8726), .ck(clk), .q(
        \pipeline/alu_out_WB [6]) );
  dp_1 \pipeline/csr/mbadaddr_reg[6]  ( .ip(n8694), .ck(clk), .q(
        \pipeline/csr/mbadaddr [6]) );
  dp_1 \pipeline/csr_rdata_WB_reg[6]  ( .ip(n8800), .ck(clk), .q(
        \pipeline/csr_rdata_WB [6]) );
  dp_1 \pipeline/store_data_WB_reg[6]  ( .ip(n8833), .ck(clk), .q(
        dmem_hwdata[6]) );
  dp_1 \pipeline/store_data_WB_reg[0]  ( .ip(n8839), .ck(clk), .q(
        dmem_hwdata[0]) );
  dp_1 \pipeline/alu_out_WB_reg[31]  ( .ip(n8701), .ck(clk), .q(
        \pipeline/alu_out_WB [31]) );
  dp_1 \pipeline/csr/mbadaddr_reg[31]  ( .ip(n8669), .ck(clk), .q(
        \pipeline/csr/mbadaddr [31]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[0]  ( .ip(n8668), .ck(clk), .q(
        htif_pcr_resp_data[0]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[1]  ( .ip(n8667), .ck(clk), .q(
        htif_pcr_resp_data[1]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[2]  ( .ip(n8666), .ck(clk), .q(
        htif_pcr_resp_data[2]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[3]  ( .ip(n8665), .ck(clk), .q(
        htif_pcr_resp_data[3]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[4]  ( .ip(n8664), .ck(clk), .q(
        htif_pcr_resp_data[4]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[5]  ( .ip(n8663), .ck(clk), .q(
        htif_pcr_resp_data[5]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[6]  ( .ip(n8662), .ck(clk), .q(
        htif_pcr_resp_data[6]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[7]  ( .ip(n8661), .ck(clk), .q(
        htif_pcr_resp_data[7]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[8]  ( .ip(n8660), .ck(clk), .q(
        htif_pcr_resp_data[8]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[9]  ( .ip(n8659), .ck(clk), .q(
        htif_pcr_resp_data[9]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[10]  ( .ip(n8658), .ck(clk), .q(
        htif_pcr_resp_data[10]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[11]  ( .ip(n8657), .ck(clk), .q(
        htif_pcr_resp_data[11]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[12]  ( .ip(n8656), .ck(clk), .q(
        htif_pcr_resp_data[12]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[13]  ( .ip(n8655), .ck(clk), .q(
        htif_pcr_resp_data[13]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[14]  ( .ip(n8654), .ck(clk), .q(
        htif_pcr_resp_data[14]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[15]  ( .ip(n8653), .ck(clk), .q(
        htif_pcr_resp_data[15]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[16]  ( .ip(n8652), .ck(clk), .q(
        htif_pcr_resp_data[16]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[17]  ( .ip(n8651), .ck(clk), .q(
        htif_pcr_resp_data[17]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[18]  ( .ip(n8650), .ck(clk), .q(
        htif_pcr_resp_data[18]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[19]  ( .ip(n8649), .ck(clk), .q(
        htif_pcr_resp_data[19]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[20]  ( .ip(n8648), .ck(clk), .q(
        htif_pcr_resp_data[20]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[21]  ( .ip(n8647), .ck(clk), .q(
        htif_pcr_resp_data[21]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[22]  ( .ip(n8646), .ck(clk), .q(
        htif_pcr_resp_data[22]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[23]  ( .ip(n8645), .ck(clk), .q(
        htif_pcr_resp_data[23]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[24]  ( .ip(n8644), .ck(clk), .q(
        htif_pcr_resp_data[24]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[25]  ( .ip(n8643), .ck(clk), .q(
        htif_pcr_resp_data[25]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[26]  ( .ip(n8642), .ck(clk), .q(
        htif_pcr_resp_data[26]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[27]  ( .ip(n8641), .ck(clk), .q(
        htif_pcr_resp_data[27]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[28]  ( .ip(n8640), .ck(clk), .q(
        htif_pcr_resp_data[28]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[29]  ( .ip(n8639), .ck(clk), .q(
        htif_pcr_resp_data[29]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[30]  ( .ip(n8638), .ck(clk), .q(
        htif_pcr_resp_data[30]) );
  dp_1 \pipeline/csr/htif_resp_data_reg[31]  ( .ip(n8637), .ck(clk), .q(
        htif_pcr_resp_data[31]) );
  dp_1 \pipeline/inst_DX_reg[14]  ( .ip(n8522), .ck(clk), .q(
        \pipeline/dmem_type[2] ) );
  dp_1 \pipeline/inst_DX_reg[26]  ( .ip(n8509), .ck(clk), .q(
        \pipeline/inst_DX [26]) );
  dp_1 \pipeline/csr/priv_stack_reg[1]  ( .ip(n10026), .ck(clk), .q(
        \pipeline/prv [0]) );
  dp_1 \pipeline/inst_DX_reg[17]  ( .ip(n8518), .ck(clk), .q(
        \pipeline/inst_DX [17]) );
  dp_1 \pipeline/csr/priv_stack_reg[2]  ( .ip(n10025), .ck(clk), .q(
        \pipeline/prv [1]) );
  dp_1 \pipeline/inst_DX_reg[27]  ( .ip(n8508), .ck(clk), .q(
        \pipeline/inst_DX [27]) );
  dp_1 \pipeline/inst_DX_reg[22]  ( .ip(n8513), .ck(clk), .q(
        \pipeline/inst_DX [22]) );
  dp_1 \pipeline/inst_DX_reg[30]  ( .ip(n8505), .ck(clk), .q(
        \pipeline/inst_DX [30]) );
  dp_1 \pipeline/inst_DX_reg[13]  ( .ip(n8523), .ck(clk), .q(dmem_hsize[1]) );
  dp_1 \pipeline/inst_DX_reg[12]  ( .ip(n8524), .ck(clk), .q(dmem_hsize[0]) );
  and2_2 U10652 ( .ip1(n14492), .ip2(n10210), .op(imem_haddr[31]) );
  inv_2 U10653 ( .ip(n16423), .op(n13552) );
  nand2_1 U10654 ( .ip1(n17387), .ip2(n10201), .op(n10700) );
  inv_1 U10655 ( .ip(n16552), .op(n10197) );
  inv_1 U10656 ( .ip(n13662), .op(n10192) );
  and2_1 U10657 ( .ip1(n10441), .ip2(n10440), .op(n10442) );
  inv_1 U10658 ( .ip(n13525), .op(n13807) );
  inv_1 U10659 ( .ip(n13727), .op(n10195) );
  inv_1 U10660 ( .ip(n17584), .op(n10194) );
  and2_1 U10661 ( .ip1(n13578), .ip2(n13895), .op(n13894) );
  inv_1 U10662 ( .ip(n13617), .op(n10188) );
  inv_1 U10663 ( .ip(n13656), .op(n10186) );
  buf_1 U10664 ( .ip(n16487), .op(n21552) );
  nor2_1 U10665 ( .ip1(\pipeline/ctrl/had_ex_WB ), .ip2(dmem_badmem_e), .op(
        n10294) );
  inv_1 U10666 ( .ip(n21082), .op(n20972) );
  nand2_1 U10667 ( .ip1(n22059), .ip2(n10201), .op(n13121) );
  inv_1 U10668 ( .ip(n13540), .op(n10185) );
  nor2_1 U10669 ( .ip1(n14289), .ip2(n14286), .op(n14287) );
  inv_1 U10670 ( .ip(n18299), .op(n14360) );
  nand2_2 U10671 ( .ip1(n16055), .ip2(n20972), .op(n10364) );
  nor2_1 U10672 ( .ip1(n22046), .ip2(n10364), .op(n17674) );
  nand2_1 U10673 ( .ip1(n14221), .ip2(n14220), .op(n14582) );
  nand2_1 U10674 ( .ip1(n14248), .ip2(n14300), .op(n14578) );
  nand2_1 U10675 ( .ip1(n17816), .ip2(n17674), .op(n17819) );
  xor2_1 U10676 ( .ip1(n10185), .ip2(n13878), .op(n10177) );
  inv_1 U10677 ( .ip(n16559), .op(n16632) );
  nand2_1 U10678 ( .ip1(n10700), .ip2(n10699), .op(n16559) );
  inv_1 U10679 ( .ip(n13022), .op(n10193) );
  inv_1 U10680 ( .ip(n13599), .op(n10191) );
  and2_1 U10681 ( .ip1(n11325), .ip2(n11324), .op(n10178) );
  and2_1 U10682 ( .ip1(ext_interrupts[19]), .ip2(\pipeline/csr/mie [27]), .op(
        n10179) );
  and2_1 U10683 ( .ip1(n11876), .ip2(n11875), .op(n10180) );
  and2_1 U10684 ( .ip1(n11600), .ip2(n11599), .op(n10181) );
  and2_1 U10685 ( .ip1(n17433), .ip2(n17431), .op(n10182) );
  inv_1 U10686 ( .ip(n13627), .op(n10189) );
  and2_1 U10687 ( .ip1(\pipeline/md/b [24]), .ip2(n15244), .op(n15245) );
  nand2_2 U10688 ( .ip1(n14545), .ip2(n10209), .op(imem_haddr[28]) );
  nand2_1 U10689 ( .ip1(n14554), .ip2(n14553), .op(n14566) );
  and2_1 U10690 ( .ip1(n14544), .ip2(n14543), .op(n10209) );
  nand2_1 U10691 ( .ip1(n14514), .ip2(n14513), .op(n14515) );
  nand2_1 U10692 ( .ip1(n14590), .ip2(n14302), .op(n14591) );
  nand2_1 U10693 ( .ip1(n14578), .ip2(n20796), .op(n14590) );
  nand2_1 U10694 ( .ip1(n14588), .ip2(n14587), .op(n20796) );
  nand2_1 U10695 ( .ip1(n14454), .ip2(n10235), .op(n14455) );
  and2_1 U10696 ( .ip1(n14507), .ip2(n14504), .op(n14508) );
  inv_1 U10697 ( .ip(n14385), .op(n14507) );
  nand2_1 U10698 ( .ip1(n20036), .ip2(n14384), .op(n14385) );
  nand2_1 U10699 ( .ip1(n17989), .ip2(n14214), .op(n14221) );
  or2_1 U10700 ( .ip1(n14555), .ip2(n14557), .op(n14565) );
  nor2_1 U10701 ( .ip1(n14585), .ip2(n14269), .op(n14270) );
  and2_1 U10702 ( .ip1(n10202), .ip2(n14531), .op(n14548) );
  and2_1 U10703 ( .ip1(n14567), .ip2(n14531), .op(n14555) );
  inv_1 U10704 ( .ip(n19489), .op(n10183) );
  nand2_1 U10705 ( .ip1(n14352), .ip2(n14353), .op(n18295) );
  nand2_1 U10706 ( .ip1(n14299), .ip2(n14301), .op(n14302) );
  nand2_1 U10707 ( .ip1(n14225), .ip2(n14303), .op(n14575) );
  and2_1 U10708 ( .ip1(n14551), .ip2(n14571), .op(n14552) );
  nand2_1 U10709 ( .ip1(n14336), .ip2(n14335), .op(n14352) );
  nand2_1 U10710 ( .ip1(n14436), .ip2(n14435), .op(n14448) );
  xnor2_1 U10711 ( .ip1(n14568), .ip2(n14567), .op(n14569) );
  xor2_2 U10712 ( .ip1(n14233), .ip2(n14234), .op(n14299) );
  and2_1 U10713 ( .ip1(n14568), .ip2(n14551), .op(n14534) );
  nand2_1 U10714 ( .ip1(n14319), .ip2(n14329), .op(n14377) );
  xor2_2 U10715 ( .ip1(n14224), .ip2(n14223), .op(n14225) );
  nand2_1 U10716 ( .ip1(n14347), .ip2(n10217), .op(n14350) );
  nand2_1 U10717 ( .ip1(n14162), .ip2(n14161), .op(n21991) );
  and2_1 U10718 ( .ip1(\pipeline/md/b [13]), .ip2(n15114), .op(n15115) );
  and2_1 U10719 ( .ip1(n14154), .ip2(n14153), .op(n14155) );
  and2_1 U10720 ( .ip1(n14326), .ip2(n14325), .op(n14327) );
  nand2_1 U10721 ( .ip1(n14328), .ip2(n14337), .op(n14331) );
  nand2_1 U10722 ( .ip1(n13579), .ip2(n13754), .op(n13752) );
  nand2_1 U10723 ( .ip1(n13749), .ip2(n10233), .op(n13750) );
  and2_1 U10724 ( .ip1(n17086), .ip2(n17085), .op(n17087) );
  and2_1 U10725 ( .ip1(n20873), .ip2(n20872), .op(n20874) );
  and2_1 U10726 ( .ip1(n17570), .ip2(n21577), .op(n17571) );
  xor2_2 U10727 ( .ip1(n17197), .ip2(n17196), .op(n17198) );
  nor2_1 U10728 ( .ip1(n13613), .ip2(n13612), .op(n13751) );
  and2_1 U10729 ( .ip1(n14035), .ip2(n14034), .op(n10238) );
  and2_1 U10730 ( .ip1(n13991), .ip2(n13909), .op(n13910) );
  and2_1 U10731 ( .ip1(n13571), .ip2(n13570), .op(n13572) );
  and2_1 U10732 ( .ip1(n17562), .ip2(n17027), .op(n17028) );
  and2_1 U10733 ( .ip1(n14241), .ip2(\pipeline/inst_DX [20]), .op(n14242) );
  and2_1 U10734 ( .ip1(n10232), .ip2(n13989), .op(n13990) );
  and2_1 U10735 ( .ip1(n13747), .ip2(n13746), .op(n13748) );
  and2_1 U10736 ( .ip1(n13872), .ip2(n13871), .op(n13873) );
  and2_1 U10737 ( .ip1(n17665), .ip2(n14032), .op(n13753) );
  and2_1 U10738 ( .ip1(n17503), .ip2(n16466), .op(n16467) );
  and2_1 U10739 ( .ip1(n17755), .ip2(n20966), .op(n17756) );
  and2_1 U10740 ( .ip1(n13782), .ip2(n13900), .op(n13783) );
  and2_1 U10741 ( .ip1(n13772), .ip2(n13861), .op(n13773) );
  and2_1 U10742 ( .ip1(n16789), .ip2(n16788), .op(n16790) );
  and2_1 U10743 ( .ip1(n13975), .ip2(n13974), .op(n13976) );
  and2_1 U10744 ( .ip1(n13800), .ip2(n17492), .op(n13801) );
  and2_1 U10745 ( .ip1(n13918), .ip2(n13917), .op(n13919) );
  and2_1 U10746 ( .ip1(n17280), .ip2(n16754), .op(n13882) );
  and2_1 U10747 ( .ip1(n16988), .ip2(n16987), .op(n16989) );
  and2_1 U10748 ( .ip1(n18930), .ip2(n19189), .op(n16610) );
  and2_1 U10749 ( .ip1(n13930), .ip2(n13929), .op(n13931) );
  and2_1 U10750 ( .ip1(n17469), .ip2(n17468), .op(n17470) );
  and2_1 U10751 ( .ip1(n13925), .ip2(n13924), .op(n13926) );
  and2_1 U10752 ( .ip1(n13933), .ip2(n13932), .op(n13934) );
  and2_1 U10753 ( .ip1(n16933), .ip2(n19051), .op(n13650) );
  and2_1 U10754 ( .ip1(n13708), .ip2(n16973), .op(n13709) );
  and2_1 U10755 ( .ip1(n17173), .ip2(n10849), .op(n13614) );
  inv_2 U10756 ( .ip(n13728), .op(n10184) );
  nor2_1 U10757 ( .ip1(n16453), .ip2(n13022), .op(n16791) );
  and2_1 U10758 ( .ip1(n17022), .ip2(n17021), .op(n17023) );
  inv_2 U10759 ( .ip(n16446), .op(n10187) );
  and2_1 U10760 ( .ip1(n10848), .ip2(n10847), .op(n10849) );
  inv_2 U10761 ( .ip(n16854), .op(n10190) );
  inv_2 U10762 ( .ip(n20903), .op(n10196) );
  nand2_2 U10763 ( .ip1(n13121), .ip2(n13120), .op(n19185) );
  mux2_1 U10764 ( .ip1(\pipeline/store_data_WB [31]), .ip2(n22069), .s(n20389), 
        .op(n8808) );
  mux2_1 U10765 ( .ip1(\pipeline/store_data_WB [29]), .ip2(n22063), .s(n17429), 
        .op(n8810) );
  inv_2 U10766 ( .ip(n10207), .op(n10198) );
  mux2_1 U10767 ( .ip1(dmem_hwdata[3]), .ip2(n22059), .s(n22067), .op(n8836)
         );
  and2_1 U10768 ( .ip1(n10895), .ip2(n10894), .op(n10896) );
  mux2_1 U10769 ( .ip1(dmem_hwdata[0]), .ip2(n22053), .s(n22067), .op(n8839)
         );
  buf_4 U10770 ( .ip(n13364), .op(n10199) );
  and2_1 U10771 ( .ip1(n13066), .ip2(n13065), .op(n17006) );
  inv_4 U10772 ( .ip(n12184), .op(n10200) );
  and2_1 U10773 ( .ip1(n10443), .ip2(n10442), .op(n10444) );
  and2_1 U10774 ( .ip1(n13521), .ip2(\pipeline/PC_DX [22]), .op(n10802) );
  inv_4 U10775 ( .ip(n12091), .op(n10201) );
  nand2_2 U10776 ( .ip1(n10289), .ip2(n10366), .op(n10454) );
  and2_1 U10777 ( .ip1(\pipeline/md/a [14]), .ip2(n20417), .op(n14648) );
  and2_1 U10778 ( .ip1(ext_interrupts[20]), .ip2(\pipeline/csr/mie [28]), .op(
        n10245) );
  and2_1 U10779 ( .ip1(n14491), .ip2(n14490), .op(n10210) );
  nor2_2 U10780 ( .ip1(n14456), .ip2(n14455), .op(n14457) );
  nand2_2 U10781 ( .ip1(n16423), .ip2(n13676), .op(n13846) );
  inv_1 U10782 ( .ip(n16690), .op(n13676) );
  nand2_2 U10783 ( .ip1(n21991), .ip2(n21992), .op(n17437) );
  nand2_2 U10784 ( .ip1(n17433), .ip2(n14439), .op(n14458) );
  nand2_4 U10785 ( .ip1(n14074), .ip2(n17669), .op(n14240) );
  nand2_2 U10786 ( .ip1(n11923), .ip2(n11922), .op(n19069) );
  nor2_4 U10787 ( .ip1(n17518), .ip2(n10239), .op(n17552) );
  nor2_1 U10788 ( .ip1(n16498), .ip2(n16626), .op(n13948) );
  nand2_1 U10789 ( .ip1(\pipeline/imm[31] ), .ip2(n14165), .op(n14337) );
  nand2_1 U10790 ( .ip1(n20035), .ip2(n20037), .op(n14445) );
  nand2_1 U10791 ( .ip1(n13678), .ip2(n20222), .op(n13863) );
  inv_1 U10792 ( .ip(n13717), .op(n13540) );
  nand2_1 U10793 ( .ip1(n12461), .ip2(n12460), .op(n16423) );
  nand2_1 U10794 ( .ip1(n20035), .ip2(n10183), .op(n14384) );
  nand2_1 U10795 ( .ip1(n14503), .ip2(n14497), .op(n14435) );
  nor2_1 U10796 ( .ip1(n13962), .ip2(n13887), .op(n12691) );
  nor2_1 U10797 ( .ip1(n10191), .ip2(n18920), .op(n11928) );
  inv_1 U10798 ( .ip(n13900), .op(n13978) );
  nor2_1 U10799 ( .ip1(n13653), .ip2(n13621), .op(n13671) );
  nor2_1 U10800 ( .ip1(n13598), .ip2(n13597), .op(n13606) );
  inv_1 U10801 ( .ip(n13746), .op(n13598) );
  nand2_1 U10802 ( .ip1(n10943), .ip2(n10942), .op(n10944) );
  nand2_1 U10803 ( .ip1(n11037), .ip2(n11036), .op(n13665) );
  nand2_1 U10804 ( .ip1(n13021), .ip2(n13020), .op(n13022) );
  and2_1 U10805 ( .ip1(n12642), .ip2(n12641), .op(n10206) );
  inv_1 U10806 ( .ip(n20222), .op(n20220) );
  nand2_1 U10807 ( .ip1(n10656), .ip2(n10655), .op(n16627) );
  and2_1 U10808 ( .ip1(n12187), .ip2(n12186), .op(n13678) );
  nand2_1 U10809 ( .ip1(n18369), .ip2(n11941), .op(n13858) );
  inv_1 U10810 ( .ip(n18369), .op(n18368) );
  inv_1 U10811 ( .ip(n13651), .op(n11941) );
  nand2_1 U10812 ( .ip1(n12885), .ip2(n12884), .op(n13878) );
  or2_1 U10813 ( .ip1(n10201), .ip2(n12883), .op(n12884) );
  nand2_1 U10814 ( .ip1(n10231), .ip2(n17297), .op(n12885) );
  inv_1 U10815 ( .ip(n12882), .op(n12883) );
  inv_1 U10816 ( .ip(n14243), .op(n14165) );
  nand2_1 U10817 ( .ip1(n14211), .ip2(n10213), .op(n14209) );
  nand2_1 U10818 ( .ip1(n14575), .ip2(n14578), .op(n14289) );
  nor4_1 U10819 ( .ip1(n17583), .ip2(n17217), .ip3(n17216), .ip4(n17215), .op(
        n17218) );
  nand2_1 U10820 ( .ip1(n12931), .ip2(n12930), .op(n12932) );
  nand2_1 U10821 ( .ip1(n22052), .ip2(n10201), .op(n12595) );
  nand2_1 U10822 ( .ip1(n12415), .ip2(n12414), .op(n16972) );
  nand2_1 U10823 ( .ip1(n12504), .ip2(n12503), .op(n16690) );
  nand4_1 U10824 ( .ip1(n16683), .ip2(n16682), .ip3(n16681), .ip4(n16680), 
        .op(n17001) );
  nand2_1 U10825 ( .ip1(n12094), .ip2(n12093), .op(n17142) );
  nand2_1 U10826 ( .ip1(n22064), .ip2(n10201), .op(n12094) );
  nand2_1 U10827 ( .ip1(n12137), .ip2(n12136), .op(n12138) );
  nand2_1 U10828 ( .ip1(n10746), .ip2(n10745), .op(n16626) );
  nand4_1 U10829 ( .ip1(n16853), .ip2(n16852), .ip3(n16851), .ip4(n21537), 
        .op(n17033) );
  and2_1 U10830 ( .ip1(n16776), .ip2(n10198), .op(n19193) );
  inv_1 U10831 ( .ip(n13878), .op(n17199) );
  nand2_1 U10832 ( .ip1(n14334), .ip2(n14331), .op(n14335) );
  nand3_1 U10833 ( .ip1(n14332), .ip2(n14333), .ip3(n14327), .op(n14336) );
  nor3_1 U10834 ( .ip1(n14448), .ip2(n14442), .ip3(n14438), .op(n14439) );
  nand2_1 U10835 ( .ip1(n14366), .ip2(n14367), .op(n14365) );
  nand2_1 U10836 ( .ip1(n14055), .ip2(n14054), .op(n14511) );
  and2_1 U10837 ( .ip1(n13977), .ip2(n13779), .op(n13904) );
  inv_1 U10838 ( .ip(n13832), .op(n13796) );
  nand2_1 U10839 ( .ip1(n13976), .ip2(n13778), .op(n13980) );
  or2_1 U10840 ( .ip1(n13771), .ip2(n14014), .op(n13774) );
  nor2_1 U10841 ( .ip1(n13766), .ip2(n13777), .op(n13775) );
  inv_1 U10842 ( .ip(n20729), .op(n13869) );
  nand2_1 U10843 ( .ip1(n11942), .ip2(n13858), .op(n11944) );
  nand2_1 U10844 ( .ip1(n11940), .ip2(n11939), .op(n11942) );
  inv_1 U10845 ( .ip(n11938), .op(n11940) );
  inv_1 U10846 ( .ip(n13770), .op(n11939) );
  nor2_1 U10847 ( .ip1(n13729), .ip2(n13726), .op(n13936) );
  nand2_1 U10848 ( .ip1(n10218), .ip2(n13725), .op(n13726) );
  nand2_1 U10849 ( .ip1(n13724), .ip2(n13723), .op(n13725) );
  nor2_1 U10850 ( .ip1(n11945), .ip2(n13981), .op(n11943) );
  nor2_1 U10851 ( .ip1(n12140), .ip2(n12139), .op(n12326) );
  nor2_1 U10852 ( .ip1(n13962), .ip2(n13889), .op(n12140) );
  nand2_1 U10853 ( .ip1(n13635), .ip2(n13634), .op(n13959) );
  nor2_1 U10854 ( .ip1(n13633), .ip2(n13632), .op(n13634) );
  nand2_1 U10855 ( .ip1(n13630), .ip2(n13629), .op(n13635) );
  nand2_1 U10856 ( .ip1(n13367), .ip2(n13366), .op(n17479) );
  nand2_1 U10857 ( .ip1(n10607), .ip2(n10606), .op(n16557) );
  nand2_1 U10858 ( .ip1(n22083), .ip2(n10201), .op(n10607) );
  nand2_1 U10859 ( .ip1(n10516), .ip2(n10515), .op(n16552) );
  nand2_1 U10860 ( .ip1(n22084), .ip2(n10201), .op(n10516) );
  nand2_1 U10861 ( .ip1(n11128), .ip2(n11127), .op(n13662) );
  nand2_1 U10862 ( .ip1(n12834), .ip2(n12833), .op(n13717) );
  nand2_1 U10863 ( .ip1(n18024), .ip2(\pipeline/PC_IF [11]), .op(n14278) );
  nand2_1 U10864 ( .ip1(\pipeline/PC_IF [14]), .ip2(n14404), .op(n14070) );
  inv_1 U10865 ( .ip(n13891), .op(n13892) );
  nand3_1 U10866 ( .ip1(n10204), .ip2(n10227), .ip3(n13890), .op(n13891) );
  nand2_1 U10867 ( .ip1(n11189), .ip2(n11188), .op(n11927) );
  nor2_1 U10868 ( .ip1(n11953), .ip2(n10216), .op(n11954) );
  nand2_1 U10869 ( .ip1(n11937), .ip2(n10230), .op(n11953) );
  nand2_1 U10870 ( .ip1(n11933), .ip2(n11932), .op(n11937) );
  nand2_1 U10871 ( .ip1(n13661), .ip2(n13660), .op(n13675) );
  nand2_1 U10872 ( .ip1(n13659), .ip2(n13658), .op(n13660) );
  nand2_1 U10873 ( .ip1(n13622), .ip2(n13671), .op(n13686) );
  nor2_1 U10874 ( .ip1(n13618), .ip2(n13908), .op(n13622) );
  nand2_1 U10875 ( .ip1(n13616), .ip2(n14002), .op(n13618) );
  nand2_1 U10876 ( .ip1(n13606), .ip2(n13605), .op(n13609) );
  nand2_1 U10877 ( .ip1(n13607), .ip2(n13606), .op(n13608) );
  inv_1 U10878 ( .ip(n13974), .op(n13607) );
  nand2_1 U10879 ( .ip1(n12741), .ip2(n12740), .op(n16445) );
  nand2_1 U10880 ( .ip1(n20221), .ip2(n20220), .op(n13862) );
  nand2_1 U10881 ( .ip1(n12231), .ip2(n12230), .op(n20222) );
  nand2_1 U10882 ( .ip1(n22062), .ip2(n10201), .op(n12231) );
  nand4_1 U10883 ( .ip1(n17454), .ip2(n17453), .ip3(n17452), .ip4(n17451), 
        .op(n20219) );
  nand2_1 U10884 ( .ip1(n12046), .ip2(n12045), .op(n19432) );
  nand2_1 U10885 ( .ip1(n22068), .ip2(n10201), .op(n12046) );
  nand2_1 U10886 ( .ip1(n13165), .ip2(n13164), .op(n13727) );
  and2_1 U10887 ( .ip1(n10790), .ip2(n10789), .op(n16498) );
  inv_1 U10888 ( .ip(n16626), .op(n13868) );
  inv_1 U10889 ( .ip(n10195), .op(n17492) );
  nand2_1 U10890 ( .ip1(n12002), .ip2(n12001), .op(n16846) );
  nand2_1 U10891 ( .ip1(n10990), .ip2(n10989), .op(n16594) );
  nand2_1 U10892 ( .ip1(n17404), .ip2(n10987), .op(n10990) );
  inv_1 U10893 ( .ip(n10944), .op(n13654) );
  nand2_2 U10894 ( .ip1(n13523), .ip2(n13522), .op(n13524) );
  nand2_1 U10895 ( .ip1(n18368), .ip2(n16914), .op(n13994) );
  nand2_1 U10896 ( .ip1(n11461), .ip2(n11460), .op(n18369) );
  inv_1 U10897 ( .ip(n11941), .op(n16914) );
  nand2_1 U10898 ( .ip1(n11370), .ip2(n11369), .op(n16935) );
  nand2_2 U10899 ( .ip1(n11279), .ip2(n11278), .op(n13601) );
  nand2_1 U10900 ( .ip1(n11416), .ip2(n11415), .op(n13651) );
  inv_1 U10901 ( .ip(n13665), .op(n11180) );
  inv_1 U10902 ( .ip(n16627), .op(n16526) );
  nand2_1 U10903 ( .ip1(n11830), .ip2(n11829), .op(n18920) );
  nand2_1 U10904 ( .ip1(n22063), .ip2(n10201), .op(n11830) );
  nor2_1 U10905 ( .ip1(n21035), .ip2(n17987), .op(n14214) );
  nand2_1 U10906 ( .ip1(n14261), .ip2(n14260), .op(n14263) );
  nand2_1 U10907 ( .ip1(n14340), .ip2(\pipeline/PC_DX [18]), .op(n14347) );
  nor2_1 U10908 ( .ip1(n14344), .ip2(n14343), .op(n14345) );
  nand2_1 U10909 ( .ip1(n14338), .ip2(n14337), .op(n14351) );
  or2_1 U10910 ( .ip1(n14445), .ip2(n14437), .op(n14442) );
  nand4_1 U10911 ( .ip1(n17206), .ip2(n17205), .ip3(n17204), .ip4(n17203), 
        .op(n21541) );
  inv_1 U10912 ( .ip(n13721), .op(n13728) );
  nand2_1 U10913 ( .ip1(n15789), .ip2(n13520), .op(n13268) );
  nand2_1 U10914 ( .ip1(n12787), .ip2(n12786), .op(n17584) );
  nand2_1 U10915 ( .ip1(n10201), .ip2(n17370), .op(n12786) );
  nor4_1 U10916 ( .ip1(n17214), .ip2(n17213), .ip3(n17212), .ip4(n17211), .op(
        n20737) );
  nand4_1 U10917 ( .ip1(n16679), .ip2(n16678), .ip3(n17527), .ip4(n18361), 
        .op(n19441) );
  nand4_1 U10918 ( .ip1(n16657), .ip2(n19187), .ip3(n18362), .ip4(n17526), 
        .op(n17520) );
  nand4_1 U10919 ( .ip1(n16660), .ip2(n16659), .ip3(n17525), .ip4(n16658), 
        .op(n20230) );
  nand4_1 U10920 ( .ip1(n19190), .ip2(n16612), .ip3(n18364), .ip4(n18929), 
        .op(n16777) );
  inv_1 U10921 ( .ip(n11508), .op(n13656) );
  nand2_1 U10922 ( .ip1(n21276), .ip2(n10201), .op(n11923) );
  nand4_1 U10923 ( .ip1(n16640), .ip2(n16639), .ip3(n16638), .ip4(n16765), 
        .op(n18944) );
  nand4_1 U10924 ( .ip1(n16631), .ip2(n16630), .ip3(n17450), .ip4(n16761), 
        .op(n18948) );
  nand2_1 U10925 ( .ip1(n11644), .ip2(n11643), .op(n17102) );
  nand2_1 U10926 ( .ip1(n22066), .ip2(n10201), .op(n11644) );
  nand2_1 U10927 ( .ip1(n22069), .ip2(n10201), .op(n11736) );
  and2_1 U10928 ( .ip1(n14194), .ip2(n14193), .op(n14210) );
  nor2_1 U10929 ( .ip1(n14192), .ip2(n14191), .op(n14193) );
  nand2_1 U10930 ( .ip1(n18024), .ip2(\pipeline/PC_IF [4]), .op(n14194) );
  inv_1 U10931 ( .ip(n14299), .op(n14248) );
  inv_1 U10932 ( .ip(n14289), .op(n14298) );
  nand2_1 U10933 ( .ip1(n14297), .ip2(n20689), .op(n14586) );
  nand2_1 U10934 ( .ip1(n14222), .ip2(n14582), .op(n14288) );
  and2_1 U10935 ( .ip1(n14305), .ip2(n14304), .op(n14306) );
  nand2_1 U10936 ( .ip1(n14589), .ip2(n14575), .op(n14305) );
  nand2_1 U10937 ( .ip1(n14079), .ip2(n14078), .op(n14363) );
  nand2_1 U10938 ( .ip1(n14077), .ip2(n14076), .op(n14079) );
  inv_1 U10939 ( .ip(n14119), .op(n14076) );
  nand2_1 U10940 ( .ip1(n18295), .ip2(n20021), .op(n14356) );
  nand4_1 U10941 ( .ip1(n10940), .ip2(n10939), .ip3(n10938), .ip4(n10937), 
        .op(n10941) );
  buf_1 U10942 ( .ip(n12683), .op(n17399) );
  nand4_1 U10943 ( .ip1(n16762), .ip2(n16761), .ip3(n16760), .ip4(n16759), 
        .op(n16772) );
  nor4_1 U10944 ( .ip1(n17221), .ip2(n17220), .ip3(n17219), .ip4(n17218), .op(
        n17241) );
  nand4_1 U10945 ( .ip1(n17462), .ip2(n16815), .ip3(n16814), .ip4(n16813), 
        .op(n16816) );
  inv_2 U10946 ( .ip(n19185), .op(n13881) );
  nand4_1 U10947 ( .ip1(n16977), .ip2(n17462), .ip3(n16976), .ip4(n16975), 
        .op(n16978) );
  nand4_1 U10948 ( .ip1(n16694), .ip2(n16693), .ip3(n16692), .ip4(n16691), 
        .op(n16695) );
  nor4_1 U10949 ( .ip1(n17052), .ip2(n17051), .ip3(n17050), .ip4(n17049), .op(
        n17152) );
  nand4_1 U10950 ( .ip1(n17148), .ip2(n17147), .ip3(n17146), .ip4(n17145), 
        .op(n17151) );
  nand4_1 U10951 ( .ip1(n16685), .ip2(n16629), .ip3(n16628), .ip4(n16658), 
        .op(n18934) );
  nand4_1 U10952 ( .ip1(n16863), .ip2(n16862), .ip3(n16861), .ip4(n16860), 
        .op(n16864) );
  nand4_1 U10953 ( .ip1(n16592), .ip2(n16686), .ip3(n16591), .ip4(n16590), 
        .op(n19426) );
  nand4_1 U10954 ( .ip1(n17284), .ip2(n17283), .ip3(n17282), .ip4(n17281), 
        .op(n17285) );
  nand4_1 U10955 ( .ip1(n16687), .ip2(n16678), .ip3(n16660), .ip4(n16587), 
        .op(n20884) );
  nand2_1 U10956 ( .ip1(n14521), .ip2(n14520), .op(n18288) );
  nand2_1 U10957 ( .ip1(n10182), .ip2(n14365), .op(n14521) );
  nand2_1 U10958 ( .ip1(n14320), .ip2(n14511), .op(n20035) );
  nor2_1 U10959 ( .ip1(n20040), .ip2(n20038), .op(n20039) );
  nand2_1 U10960 ( .ip1(n20042), .ip2(n10237), .op(n20043) );
  nand2_1 U10961 ( .ip1(n14041), .ip2(n14040), .op(n14497) );
  nor2_1 U10962 ( .ip1(n14483), .ip2(n14427), .op(n14476) );
  inv_1 U10963 ( .ip(n14528), .op(n14477) );
  or2_1 U10964 ( .ip1(n14487), .ip2(n14486), .op(n14488) );
  inv_1 U10965 ( .ip(n14485), .op(n14486) );
  nand2_1 U10966 ( .ip1(n14459), .ip2(n14528), .op(n14475) );
  nand2_1 U10967 ( .ip1(n14505), .ip2(n14506), .op(n14514) );
  nor2_1 U10968 ( .ip1(n10184), .ip2(n13881), .op(n13937) );
  nand2_1 U10969 ( .ip1(n13942), .ip2(n13941), .op(n13943) );
  nand2_1 U10970 ( .ip1(n13940), .ip2(n13939), .op(n13941) );
  inv_1 U10971 ( .ip(n13936), .op(n13942) );
  nor2_1 U10972 ( .ip1(n19193), .ip2(n13937), .op(n13940) );
  and2_1 U10973 ( .ip1(n13922), .ip2(n10225), .op(n13935) );
  nand2_1 U10974 ( .ip1(n13964), .ip2(n13963), .op(n13965) );
  inv_1 U10975 ( .ip(n13961), .op(n13964) );
  nand2_1 U10976 ( .ip1(n12596), .ip2(n16811), .op(n13922) );
  nor2_1 U10977 ( .ip1(n10193), .ip2(n13537), .op(n13538) );
  nand2_1 U10978 ( .ip1(n13656), .ip2(n18731), .op(n13770) );
  nand2_1 U10979 ( .ip1(n13722), .ip2(n13804), .op(n13723) );
  nand3_1 U10980 ( .ip1(n13863), .ip2(n13626), .ip3(n13889), .op(n13950) );
  nand2_1 U10981 ( .ip1(n13968), .ip2(n13967), .op(n13969) );
  nand3_1 U10982 ( .ip1(n13966), .ip2(n13960), .ip3(n13959), .op(n13968) );
  nand2_1 U10983 ( .ip1(n13966), .ip2(n13965), .op(n13967) );
  inv_1 U10984 ( .ip(n13958), .op(n13966) );
  nand2_1 U10985 ( .ip1(n13770), .ip2(n13858), .op(n14006) );
  nand2_1 U10986 ( .ip1(n13904), .ip2(n13903), .op(n13905) );
  nor2_1 U10987 ( .ip1(n13902), .ip2(n13901), .op(n13903) );
  nand2_1 U10988 ( .ip1(n10224), .ip2(n13861), .op(n13901) );
  nor2_1 U10989 ( .ip1(n20910), .ip2(n17177), .op(n13857) );
  inv_1 U10990 ( .ip(n17534), .op(n13856) );
  inv_1 U10991 ( .ip(n16688), .op(n13849) );
  nor2_1 U10992 ( .ip1(n17046), .ip2(n17588), .op(n13848) );
  nand2_1 U10993 ( .ip1(n10792), .ip2(n10791), .op(n10795) );
  nand3_1 U10994 ( .ip1(n13885), .ip2(n13868), .ip3(n16418), .op(n10792) );
  and2_1 U10995 ( .ip1(n16506), .ip2(n17142), .op(n13679) );
  nor2_1 U10996 ( .ip1(n13166), .ip2(n13727), .op(n13729) );
  nor2_1 U10997 ( .ip1(n13690), .ip2(n13911), .op(n13688) );
  nand2_1 U10998 ( .ip1(n13619), .ip2(n13845), .op(n13653) );
  or2_1 U10999 ( .ip1(n18368), .ip2(n13651), .op(n13619) );
  nand2_1 U11000 ( .ip1(n13628), .ip2(n13846), .op(n13629) );
  inv_1 U11001 ( .ip(n13950), .op(n13630) );
  nor2_1 U11002 ( .ip1(n13679), .ip2(n13862), .op(n13632) );
  nand4_1 U11003 ( .ip1(n12524), .ip2(n12523), .ip3(n12522), .ip4(n12521), 
        .op(n12540) );
  nand4_1 U11004 ( .ip1(n10347), .ip2(n15310), .ip3(n10330), .ip4(n17740), 
        .op(n10314) );
  nand3_1 U11005 ( .ip1(n13988), .ip2(n13987), .ip3(n13976), .op(n13989) );
  nand2_1 U11006 ( .ip1(n13776), .ip2(n13775), .op(n13785) );
  nand2_1 U11007 ( .ip1(n13774), .ip2(n13773), .op(n13776) );
  nor2_1 U11008 ( .ip1(n13869), .ip2(n16494), .op(n13876) );
  nor4_1 U11009 ( .ip1(n16598), .ip2(n16637), .ip3(n17141), .ip4(n17010), .op(
        n13890) );
  nand2_1 U11010 ( .ip1(n13865), .ip2(n13864), .op(n13866) );
  nor3_1 U11011 ( .ip1(n16900), .ip2(n13859), .ip3(n18373), .op(n13865) );
  nor4_1 U11012 ( .ip1(n17461), .ip2(n19203), .ip3(n20226), .ip4(n18924), .op(
        n13864) );
  nand2_1 U11013 ( .ip1(n13857), .ip2(n13856), .op(n13859) );
  nand2_1 U11014 ( .ip1(n13852), .ip2(n13851), .op(n13867) );
  nor4_1 U11015 ( .ip1(n16932), .ip2(n16858), .ip3(n17099), .ip4(n19438), .op(
        n13852) );
  nor2_1 U11016 ( .ip1(n13850), .ip2(n19073), .op(n13851) );
  nand2_1 U11017 ( .ip1(n13849), .ip2(n13848), .op(n13850) );
  nor2_1 U11018 ( .ip1(n11941), .ip2(n18369), .op(n11938) );
  nand2_1 U11019 ( .ip1(n12692), .ip2(n12691), .op(n13832) );
  nand2_1 U11020 ( .ip1(n11931), .ip2(n11930), .op(n11933) );
  nand2_1 U11021 ( .ip1(n11949), .ip2(n10220), .op(n11952) );
  nand2_1 U11022 ( .ip1(n11944), .ip2(n11943), .op(n11949) );
  inv_1 U11023 ( .ip(n11950), .op(n11951) );
  inv_1 U11024 ( .ip(n13917), .op(n13703) );
  or2_1 U11025 ( .ip1(n13657), .ip2(n13765), .op(n13658) );
  nor2_1 U11026 ( .ip1(n13997), .ip2(n13667), .op(n13668) );
  nor2_1 U11027 ( .ip1(n13948), .ip2(n13637), .op(n13640) );
  nand2_1 U11028 ( .ip1(n19430), .ip2(n19433), .op(n13637) );
  inv_1 U11029 ( .ip(n17006), .op(n13537) );
  xor2_1 U11030 ( .ip1(n13613), .ip2(n17006), .op(n16453) );
  nor2_1 U11031 ( .ip1(n10206), .ip2(n17457), .op(n13925) );
  nor2_1 U11032 ( .ip1(n13636), .ip2(n19432), .op(n13962) );
  nor2_1 U11033 ( .ip1(n16627), .ip2(n16632), .op(n13947) );
  nand2_1 U11034 ( .ip1(n14404), .ip2(\pipeline/PC_IF [18]), .op(n14346) );
  nand2_1 U11035 ( .ip1(n14447), .ip2(n14507), .op(n14450) );
  nand2_1 U11036 ( .ip1(n19490), .ip2(n14446), .op(n14447) );
  inv_1 U11037 ( .ip(n14445), .op(n14446) );
  nand4_1 U11038 ( .ip1(n13141), .ip2(n13140), .ip3(n13139), .ip4(n13138), 
        .op(n13157) );
  nand4_1 U11039 ( .ip1(n12908), .ip2(n12907), .ip3(n12906), .ip4(n12905), 
        .op(n12924) );
  nand4_1 U11040 ( .ip1(n12863), .ip2(n12862), .ip3(n12861), .ip4(n12860), 
        .op(n12874) );
  nand4_1 U11041 ( .ip1(n12998), .ip2(n12997), .ip3(n12996), .ip4(n12995), 
        .op(n13014) );
  nand4_1 U11042 ( .ip1(n12619), .ip2(n12618), .ip3(n12617), .ip4(n12616), 
        .op(n12635) );
  nand4_1 U11043 ( .ip1(n12510), .ip2(n12509), .ip3(n12508), .ip4(n12507), 
        .op(n12511) );
  nor4_1 U11044 ( .ip1(n12540), .ip2(n12539), .ip3(n12538), .ip4(n12537), .op(
        n12541) );
  nand4_1 U11045 ( .ip1(n12532), .ip2(n12531), .ip3(n12530), .ip4(n12529), 
        .op(n12538) );
  nand4_1 U11046 ( .ip1(n12536), .ip2(n12535), .ip3(n12534), .ip4(n12533), 
        .op(n12537) );
  nand4_1 U11047 ( .ip1(n12528), .ip2(n12527), .ip3(n12526), .ip4(n12525), 
        .op(n12539) );
  nor4_1 U11048 ( .ip1(n10436), .ip2(n10435), .ip3(n10434), .ip4(n10451), .op(
        n10439) );
  nand4_1 U11049 ( .ip1(n13343), .ip2(n13342), .ip3(n13341), .ip4(n13340), 
        .op(n13359) );
  nand4_1 U11050 ( .ip1(n13243), .ip2(n13242), .ip3(n13241), .ip4(n13240), 
        .op(n13259) );
  nand4_1 U11051 ( .ip1(n12114), .ip2(n12113), .ip3(n12112), .ip4(n12111), 
        .op(n12130) );
  nand4_1 U11052 ( .ip1(n12811), .ip2(n12810), .ip3(n12809), .ip4(n12808), 
        .op(n12827) );
  nand4_1 U11053 ( .ip1(n10403), .ip2(n10402), .ip3(n10401), .ip4(n10400), 
        .op(n10429) );
  nand4_1 U11054 ( .ip1(n11393), .ip2(n11392), .ip3(n11391), .ip4(n11390), 
        .op(n11409) );
  nand4_1 U11055 ( .ip1(n11152), .ip2(n11151), .ip3(n11150), .ip4(n11149), 
        .op(n11163) );
  nand4_1 U11056 ( .ip1(n10968), .ip2(n10967), .ip3(n10966), .ip4(n10965), 
        .op(n10979) );
  nand4_1 U11057 ( .ip1(n11440), .ip2(n11439), .ip3(n11438), .ip4(n11437), 
        .op(n11451) );
  nand4_1 U11058 ( .ip1(n12254), .ip2(n12253), .ip3(n12252), .ip4(n12251), 
        .op(n12270) );
  nand4_1 U11059 ( .ip1(n10920), .ip2(n10919), .ip3(n10918), .ip4(n10917), 
        .op(n10936) );
  nand4_1 U11060 ( .ip1(n11105), .ip2(n11104), .ip3(n11103), .ip4(n11102), 
        .op(n11121) );
  nand4_1 U11061 ( .ip1(n10822), .ip2(n10821), .ip3(n10820), .ip4(n10819), 
        .op(n10838) );
  nand4_1 U11062 ( .ip1(n10826), .ip2(n10825), .ip3(n10824), .ip4(n10823), 
        .op(n10837) );
  nand4_1 U11063 ( .ip1(n10834), .ip2(n10833), .ip3(n10832), .ip4(n10831), 
        .op(n10835) );
  nand4_1 U11064 ( .ip1(n10830), .ip2(n10829), .ip3(n10828), .ip4(n10827), 
        .op(n10836) );
  nand4_1 U11065 ( .ip1(n10808), .ip2(n10807), .ip3(n10806), .ip4(n10805), 
        .op(n10809) );
  nand4_1 U11066 ( .ip1(n11011), .ip2(n11010), .ip3(n11009), .ip4(n11008), 
        .op(n11027) );
  nand4_1 U11067 ( .ip1(n11259), .ip2(n11258), .ip3(n11257), .ip4(n11256), 
        .op(n11270) );
  nand4_1 U11068 ( .ip1(n11212), .ip2(n11211), .ip3(n11210), .ip4(n11209), 
        .op(n11228) );
  nand4_1 U11069 ( .ip1(n12438), .ip2(n12437), .ip3(n12436), .ip4(n12435), 
        .op(n12454) );
  nand4_1 U11070 ( .ip1(n12349), .ip2(n12348), .ip3(n12347), .ip4(n12346), 
        .op(n12365) );
  nand4_1 U11071 ( .ip1(n11853), .ip2(n11852), .ip3(n11851), .ip4(n11850), 
        .op(n11869) );
  nand4_1 U11072 ( .ip1(n11978), .ip2(n11977), .ip3(n11976), .ip4(n11975), 
        .op(n11994) );
  nand4_1 U11073 ( .ip1(n10723), .ip2(n10722), .ip3(n10721), .ip4(n10720), 
        .op(n10739) );
  nand4_1 U11074 ( .ip1(n11577), .ip2(n11576), .ip3(n11575), .ip4(n11574), 
        .op(n11593) );
  inv_1 U11075 ( .ip(n13524), .op(n13870) );
  inv_1 U11076 ( .ip(n17479), .op(n16608) );
  xor2_1 U11077 ( .ip1(n17199), .ip2(n16913), .op(n16443) );
  nand2_1 U11078 ( .ip1(n17040), .ip2(n17042), .op(n13930) );
  nor2_1 U11079 ( .ip1(n16506), .ip2(n17142), .op(n13887) );
  nand2_1 U11080 ( .ip1(n17142), .ip2(n16506), .op(n13889) );
  inv_1 U11081 ( .ip(n12138), .op(n16506) );
  inv_1 U11082 ( .ip(n19432), .op(n19430) );
  inv_1 U11083 ( .ip(n10206), .op(n17456) );
  inv_1 U11084 ( .ip(n16846), .op(n13636) );
  nand2_1 U11085 ( .ip1(n10197), .ip2(n13666), .op(n13997) );
  nand2_1 U11086 ( .ip1(n16593), .ip2(n10944), .op(n13993) );
  inv_1 U11087 ( .ip(n16594), .op(n16593) );
  nand4_1 U11088 ( .ip1(n16649), .ip2(n19188), .ip3(n18363), .ip4(n18932), 
        .op(n17519) );
  and2_1 U11089 ( .ip1(n13223), .ip2(n13222), .op(n10207) );
  nor4_1 U11090 ( .ip1(n16946), .ip2(n16945), .ip3(n16944), .ip4(n16943), .op(
        n17106) );
  nand2_1 U11091 ( .ip1(n17073), .ip2(n17100), .op(n13974) );
  inv_1 U11092 ( .ip(n17102), .op(n17100) );
  nand2_1 U11093 ( .ip1(n11934), .ip2(n10196), .op(n13900) );
  nand4_1 U11094 ( .ip1(n13486), .ip2(n13485), .ip3(n13484), .ip4(n13483), 
        .op(n13514) );
  nor2_1 U11095 ( .ip1(n14280), .ip2(n14279), .op(n14281) );
  nand2_1 U11096 ( .ip1(n14278), .ip2(n14277), .op(n14279) );
  nor2_1 U11097 ( .ip1(n14275), .ip2(n14276), .op(n14280) );
  and2_1 U11098 ( .ip1(n14071), .ip2(n14070), .op(n14072) );
  nand2_1 U11099 ( .ip1(n14399), .ip2(\pipeline/PC_DX [14]), .op(n14073) );
  nor2_1 U11100 ( .ip1(n14069), .ip2(n14068), .op(n14071) );
  nand2_1 U11101 ( .ip1(n14114), .ip2(n14113), .op(n14118) );
  nand2_1 U11102 ( .ip1(\pipeline/PC_DX [15]), .ip2(n14399), .op(n14114) );
  nand2_1 U11103 ( .ip1(n14413), .ip2(\pipeline/PC_DX [19]), .op(n14332) );
  nand2_1 U11104 ( .ip1(n14089), .ip2(n14337), .op(n14349) );
  nand4_1 U11105 ( .ip1(n17431), .ip2(n14440), .ip3(n18285), .ip4(n14365), 
        .op(n14438) );
  or2_1 U11106 ( .ip1(n14517), .ip2(n14448), .op(n14441) );
  nand4_1 U11107 ( .ip1(n12073), .ip2(n12072), .ip3(n12071), .ip4(n12070), 
        .op(n12084) );
  nand4_1 U11108 ( .ip1(n10680), .ip2(n10679), .ip3(n10678), .ip4(n10677), 
        .op(n10691) );
  nand4_1 U11109 ( .ip1(n12211), .ip2(n12210), .ip3(n12209), .ip4(n12208), 
        .op(n12222) );
  nand4_1 U11110 ( .ip1(n12301), .ip2(n12300), .ip3(n12299), .ip4(n12298), 
        .op(n12312) );
  nand4_1 U11111 ( .ip1(n11349), .ip2(n11348), .ip3(n11347), .ip4(n11346), 
        .op(n11360) );
  nand4_1 U11112 ( .ip1(n11808), .ip2(n11807), .ip3(n11806), .ip4(n11805), 
        .op(n11819) );
  nand4_1 U11113 ( .ip1(n11624), .ip2(n11623), .ip3(n11622), .ip4(n11621), 
        .op(n11635) );
  nand4_1 U11114 ( .ip1(n13127), .ip2(n13126), .ip3(n13125), .ip4(n13124), 
        .op(n13128) );
  nor4_1 U11115 ( .ip1(n13157), .ip2(n13156), .ip3(n13155), .ip4(n13154), .op(
        n13158) );
  nand4_1 U11116 ( .ip1(n13149), .ip2(n13148), .ip3(n13147), .ip4(n13146), 
        .op(n13155) );
  nand4_1 U11117 ( .ip1(n13153), .ip2(n13152), .ip3(n13151), .ip4(n13150), 
        .op(n13154) );
  nand4_1 U11118 ( .ip1(n13145), .ip2(n13144), .ip3(n13143), .ip4(n13142), 
        .op(n13156) );
  nand4_1 U11119 ( .ip1(n12894), .ip2(n12893), .ip3(n12892), .ip4(n12891), 
        .op(n12895) );
  nor4_1 U11120 ( .ip1(n12924), .ip2(n12923), .ip3(n12922), .ip4(n12921), .op(
        n12925) );
  nand4_1 U11121 ( .ip1(n12916), .ip2(n12915), .ip3(n12914), .ip4(n12913), 
        .op(n12922) );
  nand4_1 U11122 ( .ip1(n12920), .ip2(n12919), .ip3(n12918), .ip4(n12917), 
        .op(n12921) );
  nand4_1 U11123 ( .ip1(n12912), .ip2(n12911), .ip3(n12910), .ip4(n12909), 
        .op(n12923) );
  nand4_1 U11124 ( .ip1(n13416), .ip2(n13415), .ip3(n13414), .ip4(n13413), 
        .op(n13435) );
  nand4_1 U11125 ( .ip1(n13298), .ip2(n13297), .ip3(n13296), .ip4(n13295), 
        .op(n13309) );
  nand4_1 U11126 ( .ip1(n13198), .ip2(n13197), .ip3(n13196), .ip4(n13195), 
        .op(n13199) );
  nand4_1 U11127 ( .ip1(n13194), .ip2(n13193), .ip3(n13192), .ip4(n13191), 
        .op(n13200) );
  nand4_1 U11128 ( .ip1(n13186), .ip2(n13185), .ip3(n13184), .ip4(n13183), 
        .op(n13202) );
  nand4_1 U11129 ( .ip1(n13190), .ip2(n13189), .ip3(n13188), .ip4(n13187), 
        .op(n13201) );
  nand4_1 U11130 ( .ip1(n13174), .ip2(n13173), .ip3(n13172), .ip4(n13171), 
        .op(n13206) );
  nand4_1 U11131 ( .ip1(n13096), .ip2(n13095), .ip3(n13094), .ip4(n13093), 
        .op(n13107) );
  nand4_1 U11132 ( .ip1(n12845), .ip2(n12844), .ip3(n12843), .ip4(n12842), 
        .op(n12846) );
  nor4_1 U11133 ( .ip1(n12875), .ip2(n12874), .ip3(n12873), .ip4(n12872), .op(
        n12876) );
  nand4_1 U11134 ( .ip1(n12867), .ip2(n12866), .ip3(n12865), .ip4(n12864), 
        .op(n12873) );
  nand4_1 U11135 ( .ip1(n12859), .ip2(n12858), .ip3(n12857), .ip4(n12856), 
        .op(n12875) );
  nand4_1 U11136 ( .ip1(n12871), .ip2(n12870), .ip3(n12869), .ip4(n12868), 
        .op(n12872) );
  nand4_1 U11137 ( .ip1(n12766), .ip2(n12765), .ip3(n12764), .ip4(n12763), 
        .op(n12777) );
  nand4_1 U11138 ( .ip1(n12956), .ip2(n12955), .ip3(n12954), .ip4(n12953), 
        .op(n12967) );
  nand4_1 U11139 ( .ip1(n12984), .ip2(n12983), .ip3(n12982), .ip4(n12981), 
        .op(n12985) );
  nor4_1 U11140 ( .ip1(n13014), .ip2(n13013), .ip3(n13012), .ip4(n13011), .op(
        n13015) );
  nand4_1 U11141 ( .ip1(n13006), .ip2(n13005), .ip3(n13004), .ip4(n13003), 
        .op(n13012) );
  nand4_1 U11142 ( .ip1(n13010), .ip2(n13009), .ip3(n13008), .ip4(n13007), 
        .op(n13011) );
  nand4_1 U11143 ( .ip1(n13002), .ip2(n13001), .ip3(n13000), .ip4(n12999), 
        .op(n13013) );
  nand4_1 U11144 ( .ip1(n13046), .ip2(n13045), .ip3(n13044), .ip4(n13043), 
        .op(n13057) );
  nand4_1 U11145 ( .ip1(n12605), .ip2(n12604), .ip3(n12603), .ip4(n12602), 
        .op(n12606) );
  nor4_1 U11146 ( .ip1(n12635), .ip2(n12634), .ip3(n12633), .ip4(n12632), .op(
        n12636) );
  nand4_1 U11147 ( .ip1(n12627), .ip2(n12626), .ip3(n12625), .ip4(n12624), 
        .op(n12633) );
  nand4_1 U11148 ( .ip1(n12631), .ip2(n12630), .ip3(n12629), .ip4(n12628), 
        .op(n12632) );
  nand4_1 U11149 ( .ip1(n12623), .ip2(n12622), .ip3(n12621), .ip4(n12620), 
        .op(n12634) );
  nand4_1 U11150 ( .ip1(n12575), .ip2(n12574), .ip3(n12573), .ip4(n12572), 
        .op(n12586) );
  nand4_1 U11151 ( .ip1(n12666), .ip2(n12665), .ip3(n12664), .ip4(n12663), 
        .op(n12677) );
  nand4_1 U11152 ( .ip1(n12716), .ip2(n12715), .ip3(n12714), .ip4(n12713), 
        .op(n12732) );
  nand4_1 U11153 ( .ip1(n13329), .ip2(n13328), .ip3(n13327), .ip4(n13326), 
        .op(n13330) );
  nor4_1 U11154 ( .ip1(n13359), .ip2(n13358), .ip3(n13357), .ip4(n13356), .op(
        n13360) );
  nand4_1 U11155 ( .ip1(n13351), .ip2(n13350), .ip3(n13349), .ip4(n13348), 
        .op(n13357) );
  nand4_1 U11156 ( .ip1(n13355), .ip2(n13354), .ip3(n13353), .ip4(n13352), 
        .op(n13356) );
  nand4_1 U11157 ( .ip1(n13347), .ip2(n13346), .ip3(n13345), .ip4(n13344), 
        .op(n13358) );
  nand4_1 U11158 ( .ip1(n13229), .ip2(n13228), .ip3(n13227), .ip4(n13226), 
        .op(n13230) );
  nor4_1 U11159 ( .ip1(n13259), .ip2(n13258), .ip3(n13257), .ip4(n13256), .op(
        n13260) );
  nand4_1 U11160 ( .ip1(n13251), .ip2(n13250), .ip3(n13249), .ip4(n13248), 
        .op(n13257) );
  nand4_1 U11161 ( .ip1(n13255), .ip2(n13254), .ip3(n13253), .ip4(n13252), 
        .op(n13256) );
  nand4_1 U11162 ( .ip1(n13247), .ip2(n13246), .ip3(n13245), .ip4(n13244), 
        .op(n13258) );
  nand4_1 U11163 ( .ip1(n12396), .ip2(n12395), .ip3(n12394), .ip4(n12393), 
        .op(n12407) );
  nand4_1 U11164 ( .ip1(n12485), .ip2(n12484), .ip3(n12483), .ip4(n12482), 
        .op(n12496) );
  nand4_1 U11165 ( .ip1(n12026), .ip2(n12025), .ip3(n12024), .ip4(n12023), 
        .op(n12037) );
  nand4_1 U11166 ( .ip1(n12100), .ip2(n12099), .ip3(n12098), .ip4(n12097), 
        .op(n12101) );
  nor4_1 U11167 ( .ip1(n12130), .ip2(n12129), .ip3(n12128), .ip4(n12127), .op(
        n12131) );
  nand4_1 U11168 ( .ip1(n12122), .ip2(n12121), .ip3(n12120), .ip4(n12119), 
        .op(n12128) );
  nand4_1 U11169 ( .ip1(n12126), .ip2(n12125), .ip3(n12124), .ip4(n12123), 
        .op(n12127) );
  nand4_1 U11170 ( .ip1(n12118), .ip2(n12117), .ip3(n12116), .ip4(n12115), 
        .op(n12129) );
  nand4_1 U11171 ( .ip1(n12797), .ip2(n12796), .ip3(n12795), .ip4(n12794), 
        .op(n12798) );
  nor4_1 U11172 ( .ip1(n12827), .ip2(n12826), .ip3(n12825), .ip4(n12824), .op(
        n12828) );
  nand4_1 U11173 ( .ip1(n12819), .ip2(n12818), .ip3(n12817), .ip4(n12816), 
        .op(n12825) );
  nand4_1 U11174 ( .ip1(n12823), .ip2(n12822), .ip3(n12821), .ip4(n12820), 
        .op(n12824) );
  nand4_1 U11175 ( .ip1(n12815), .ip2(n12814), .ip3(n12813), .ip4(n12812), 
        .op(n12826) );
  nand4_1 U11176 ( .ip1(n10385), .ip2(n10384), .ip3(n10383), .ip4(n10382), 
        .op(n10386) );
  nor4_1 U11177 ( .ip1(n10429), .ip2(n10428), .ip3(n10427), .ip4(n10426), .op(
        n10430) );
  nand4_1 U11178 ( .ip1(n10416), .ip2(n10415), .ip3(n10414), .ip4(n10413), 
        .op(n10427) );
  nand4_1 U11179 ( .ip1(n10425), .ip2(n10424), .ip3(n10423), .ip4(n10422), 
        .op(n10426) );
  nand4_1 U11180 ( .ip1(n10409), .ip2(n10408), .ip3(n10407), .ip4(n10406), 
        .op(n10428) );
  nand4_1 U11181 ( .ip1(n10771), .ip2(n10770), .ip3(n10769), .ip4(n10768), 
        .op(n10782) );
  nand4_1 U11182 ( .ip1(n10587), .ip2(n10586), .ip3(n10585), .ip4(n10584), 
        .op(n10598) );
  nand4_1 U11183 ( .ip1(n10485), .ip2(n10484), .ip3(n10483), .ip4(n10482), 
        .op(n10502) );
  nand4_1 U11184 ( .ip1(n10540), .ip2(n10539), .ip3(n10538), .ip4(n10537), 
        .op(n10556) );
  nand4_1 U11185 ( .ip1(n11379), .ip2(n11378), .ip3(n11377), .ip4(n11376), 
        .op(n11380) );
  nor4_1 U11186 ( .ip1(n11409), .ip2(n11408), .ip3(n11407), .ip4(n11406), .op(
        n11410) );
  nand4_1 U11187 ( .ip1(n11401), .ip2(n11400), .ip3(n11399), .ip4(n11398), 
        .op(n11407) );
  nand4_1 U11188 ( .ip1(n11405), .ip2(n11404), .ip3(n11403), .ip4(n11402), 
        .op(n11406) );
  nand4_1 U11189 ( .ip1(n11397), .ip2(n11396), .ip3(n11395), .ip4(n11394), 
        .op(n11408) );
  nand4_1 U11190 ( .ip1(n11061), .ip2(n11060), .ip3(n11059), .ip4(n11058), 
        .op(n11072) );
  nand4_1 U11191 ( .ip1(n11134), .ip2(n11133), .ip3(n11132), .ip4(n11131), 
        .op(n11135) );
  nor4_1 U11192 ( .ip1(n11164), .ip2(n11163), .ip3(n11162), .ip4(n11161), .op(
        n11165) );
  nand4_1 U11193 ( .ip1(n11156), .ip2(n11155), .ip3(n11154), .ip4(n11153), 
        .op(n11162) );
  nand4_1 U11194 ( .ip1(n11148), .ip2(n11147), .ip3(n11146), .ip4(n11145), 
        .op(n11164) );
  nand4_1 U11195 ( .ip1(n11160), .ip2(n11159), .ip3(n11158), .ip4(n11157), 
        .op(n11161) );
  nand4_1 U11196 ( .ip1(n10875), .ip2(n10874), .ip3(n10873), .ip4(n10872), 
        .op(n10886) );
  nand4_1 U11197 ( .ip1(n10883), .ip2(n10882), .ip3(n10881), .ip4(n10880), 
        .op(n10884) );
  nand4_1 U11198 ( .ip1(n10871), .ip2(n10870), .ip3(n10869), .ip4(n10868), 
        .op(n10887) );
  nand4_1 U11199 ( .ip1(n10879), .ip2(n10878), .ip3(n10877), .ip4(n10876), 
        .op(n10885) );
  nand4_1 U11200 ( .ip1(n10857), .ip2(n10856), .ip3(n10855), .ip4(n10854), 
        .op(n10858) );
  nand4_1 U11201 ( .ip1(n10950), .ip2(n10949), .ip3(n10948), .ip4(n10947), 
        .op(n10951) );
  nor4_1 U11202 ( .ip1(n10980), .ip2(n10979), .ip3(n10978), .ip4(n10977), .op(
        n10981) );
  nand4_1 U11203 ( .ip1(n10972), .ip2(n10971), .ip3(n10970), .ip4(n10969), 
        .op(n10978) );
  nand4_1 U11204 ( .ip1(n10964), .ip2(n10963), .ip3(n10962), .ip4(n10961), 
        .op(n10980) );
  nand4_1 U11205 ( .ip1(n10976), .ip2(n10975), .ip3(n10974), .ip4(n10973), 
        .op(n10977) );
  nand4_1 U11206 ( .ip1(n11532), .ip2(n11531), .ip3(n11530), .ip4(n11529), 
        .op(n11543) );
  nand4_1 U11207 ( .ip1(n11422), .ip2(n11421), .ip3(n11420), .ip4(n11419), 
        .op(n11423) );
  nor4_1 U11208 ( .ip1(n11452), .ip2(n11451), .ip3(n11450), .ip4(n11449), .op(
        n11453) );
  nand4_1 U11209 ( .ip1(n11444), .ip2(n11443), .ip3(n11442), .ip4(n11441), 
        .op(n11450) );
  nand4_1 U11210 ( .ip1(n11436), .ip2(n11435), .ip3(n11434), .ip4(n11433), 
        .op(n11452) );
  nand4_1 U11211 ( .ip1(n11448), .ip2(n11447), .ip3(n11446), .ip4(n11445), 
        .op(n11449) );
  nand4_1 U11212 ( .ip1(n10633), .ip2(n10632), .ip3(n10631), .ip4(n10630), 
        .op(n10649) );
  nand4_1 U11213 ( .ip1(n12163), .ip2(n12162), .ip3(n12161), .ip4(n12160), 
        .op(n12179) );
  nand4_1 U11214 ( .ip1(n12240), .ip2(n12239), .ip3(n12238), .ip4(n12237), 
        .op(n12241) );
  nor4_1 U11215 ( .ip1(n12270), .ip2(n12269), .ip3(n12268), .ip4(n12267), .op(
        n12271) );
  nand4_1 U11216 ( .ip1(n12262), .ip2(n12261), .ip3(n12260), .ip4(n12259), 
        .op(n12268) );
  nand4_1 U11217 ( .ip1(n12266), .ip2(n12265), .ip3(n12264), .ip4(n12263), 
        .op(n12267) );
  nand4_1 U11218 ( .ip1(n12258), .ip2(n12257), .ip3(n12256), .ip4(n12255), 
        .op(n12269) );
  nand4_1 U11219 ( .ip1(n10906), .ip2(n10905), .ip3(n10904), .ip4(n10903), 
        .op(n10907) );
  nor4_1 U11220 ( .ip1(n10936), .ip2(n10935), .ip3(n10934), .ip4(n10933), .op(
        n10937) );
  nand4_1 U11221 ( .ip1(n10928), .ip2(n10927), .ip3(n10926), .ip4(n10925), 
        .op(n10934) );
  nand4_1 U11222 ( .ip1(n10932), .ip2(n10931), .ip3(n10930), .ip4(n10929), 
        .op(n10933) );
  nand4_1 U11223 ( .ip1(n10924), .ip2(n10923), .ip3(n10922), .ip4(n10921), 
        .op(n10935) );
  nand4_1 U11224 ( .ip1(n11091), .ip2(n11090), .ip3(n11089), .ip4(n11088), 
        .op(n11092) );
  nor4_1 U11225 ( .ip1(n11121), .ip2(n11120), .ip3(n11119), .ip4(n11118), .op(
        n11122) );
  nand4_1 U11226 ( .ip1(n11113), .ip2(n11112), .ip3(n11111), .ip4(n11110), 
        .op(n11119) );
  nand4_1 U11227 ( .ip1(n11117), .ip2(n11116), .ip3(n11115), .ip4(n11114), 
        .op(n11118) );
  nand4_1 U11228 ( .ip1(n11109), .ip2(n11108), .ip3(n11107), .ip4(n11106), 
        .op(n11120) );
  nand4_1 U11229 ( .ip1(n10842), .ip2(n10841), .ip3(n10840), .ip4(n10839), 
        .op(n14056) );
  nor4_1 U11230 ( .ip1(n10838), .ip2(n10837), .ip3(n10836), .ip4(n10835), .op(
        n10839) );
  nand4_1 U11231 ( .ip1(n10997), .ip2(n10996), .ip3(n10995), .ip4(n10994), 
        .op(n10998) );
  nor4_1 U11232 ( .ip1(n11027), .ip2(n11026), .ip3(n11025), .ip4(n11024), .op(
        n11028) );
  nand4_1 U11233 ( .ip1(n11019), .ip2(n11018), .ip3(n11017), .ip4(n11016), 
        .op(n11025) );
  nand4_1 U11234 ( .ip1(n11023), .ip2(n11022), .ip3(n11021), .ip4(n11020), 
        .op(n11024) );
  nand4_1 U11235 ( .ip1(n11015), .ip2(n11014), .ip3(n11013), .ip4(n11012), 
        .op(n11026) );
  nand4_1 U11236 ( .ip1(n11302), .ip2(n11301), .ip3(n11300), .ip4(n11299), 
        .op(n11318) );
  nand4_1 U11237 ( .ip1(n11760), .ip2(n11759), .ip3(n11758), .ip4(n11757), 
        .op(n11776) );
  nand4_1 U11238 ( .ip1(n11241), .ip2(n11240), .ip3(n11239), .ip4(n11238), 
        .op(n11242) );
  nor4_1 U11239 ( .ip1(n11271), .ip2(n11270), .ip3(n11269), .ip4(n11268), .op(
        n11272) );
  nand4_1 U11240 ( .ip1(n11263), .ip2(n11262), .ip3(n11261), .ip4(n11260), 
        .op(n11269) );
  nand4_1 U11241 ( .ip1(n11255), .ip2(n11254), .ip3(n11253), .ip4(n11252), 
        .op(n11271) );
  nand4_1 U11242 ( .ip1(n11267), .ip2(n11266), .ip3(n11265), .ip4(n11264), 
        .op(n11268) );
  nand4_1 U11243 ( .ip1(n11901), .ip2(n11900), .ip3(n11899), .ip4(n11898), 
        .op(n11912) );
  nand4_1 U11244 ( .ip1(n11909), .ip2(n11908), .ip3(n11907), .ip4(n11906), 
        .op(n11910) );
  nand4_1 U11245 ( .ip1(n11897), .ip2(n11896), .ip3(n11895), .ip4(n11894), 
        .op(n11913) );
  nand4_1 U11246 ( .ip1(n11905), .ip2(n11904), .ip3(n11903), .ip4(n11902), 
        .op(n11911) );
  nand4_1 U11247 ( .ip1(n11883), .ip2(n11882), .ip3(n11881), .ip4(n11880), 
        .op(n11884) );
  nand4_1 U11248 ( .ip1(n11198), .ip2(n11197), .ip3(n11196), .ip4(n11195), 
        .op(n11199) );
  nor4_1 U11249 ( .ip1(n11228), .ip2(n11227), .ip3(n11226), .ip4(n11225), .op(
        n11229) );
  nand4_1 U11250 ( .ip1(n11220), .ip2(n11219), .ip3(n11218), .ip4(n11217), 
        .op(n11226) );
  nand4_1 U11251 ( .ip1(n11224), .ip2(n11223), .ip3(n11222), .ip4(n11221), 
        .op(n11225) );
  nand4_1 U11252 ( .ip1(n11216), .ip2(n11215), .ip3(n11214), .ip4(n11213), 
        .op(n11227) );
  nand4_1 U11253 ( .ip1(n12424), .ip2(n12423), .ip3(n12422), .ip4(n12421), 
        .op(n12425) );
  nor4_1 U11254 ( .ip1(n12454), .ip2(n12453), .ip3(n12452), .ip4(n12451), .op(
        n12455) );
  nand4_1 U11255 ( .ip1(n12446), .ip2(n12445), .ip3(n12444), .ip4(n12443), 
        .op(n12452) );
  nand4_1 U11256 ( .ip1(n12450), .ip2(n12449), .ip3(n12448), .ip4(n12447), 
        .op(n12451) );
  nand4_1 U11257 ( .ip1(n12442), .ip2(n12441), .ip3(n12440), .ip4(n12439), 
        .op(n12453) );
  nand4_1 U11258 ( .ip1(n12335), .ip2(n12334), .ip3(n12333), .ip4(n12332), 
        .op(n12336) );
  nor4_1 U11259 ( .ip1(n12365), .ip2(n12364), .ip3(n12363), .ip4(n12362), .op(
        n12366) );
  nand4_1 U11260 ( .ip1(n12357), .ip2(n12356), .ip3(n12355), .ip4(n12354), 
        .op(n12363) );
  nand4_1 U11261 ( .ip1(n12361), .ip2(n12360), .ip3(n12359), .ip4(n12358), 
        .op(n12362) );
  nand4_1 U11262 ( .ip1(n12353), .ip2(n12352), .ip3(n12351), .ip4(n12350), 
        .op(n12364) );
  nand4_1 U11263 ( .ip1(n11839), .ip2(n11838), .ip3(n11837), .ip4(n11836), 
        .op(n11840) );
  nor4_1 U11264 ( .ip1(n11869), .ip2(n11868), .ip3(n11867), .ip4(n11866), .op(
        n11870) );
  nand4_1 U11265 ( .ip1(n11861), .ip2(n11860), .ip3(n11859), .ip4(n11858), 
        .op(n11867) );
  nand4_1 U11266 ( .ip1(n11865), .ip2(n11864), .ip3(n11863), .ip4(n11862), 
        .op(n11866) );
  nand4_1 U11267 ( .ip1(n11857), .ip2(n11856), .ip3(n11855), .ip4(n11854), 
        .op(n11868) );
  nand4_1 U11268 ( .ip1(n11484), .ip2(n11483), .ip3(n11482), .ip4(n11481), 
        .op(n11500) );
  nand4_1 U11269 ( .ip1(n11964), .ip2(n11963), .ip3(n11962), .ip4(n11961), 
        .op(n11965) );
  nor4_1 U11270 ( .ip1(n11994), .ip2(n11993), .ip3(n11992), .ip4(n11991), .op(
        n11995) );
  nand4_1 U11271 ( .ip1(n11986), .ip2(n11985), .ip3(n11984), .ip4(n11983), 
        .op(n11992) );
  nand4_1 U11272 ( .ip1(n11990), .ip2(n11989), .ip3(n11988), .ip4(n11987), 
        .op(n11991) );
  nand4_1 U11273 ( .ip1(n11982), .ip2(n11981), .ip3(n11980), .ip4(n11979), 
        .op(n11993) );
  nand4_1 U11274 ( .ip1(n10709), .ip2(n10708), .ip3(n10707), .ip4(n10706), 
        .op(n10710) );
  nor4_1 U11275 ( .ip1(n10739), .ip2(n10738), .ip3(n10737), .ip4(n10736), .op(
        n10740) );
  nand4_1 U11276 ( .ip1(n10731), .ip2(n10730), .ip3(n10729), .ip4(n10728), 
        .op(n10737) );
  nand4_1 U11277 ( .ip1(n10735), .ip2(n10734), .ip3(n10733), .ip4(n10732), 
        .op(n10736) );
  nand4_1 U11278 ( .ip1(n10727), .ip2(n10726), .ip3(n10725), .ip4(n10724), 
        .op(n10738) );
  nor4_1 U11279 ( .ip1(n10298), .ip2(n10436), .ip3(n10435), .ip4(n10297), .op(
        n10312) );
  nand4_1 U11280 ( .ip1(n11715), .ip2(n11714), .ip3(n11713), .ip4(n11712), 
        .op(n11726) );
  nand2_1 U11281 ( .ip1(n16496), .ip2(n13843), .op(n14024) );
  nand4_1 U11282 ( .ip1(n11667), .ip2(n11666), .ip3(n11665), .ip4(n11664), 
        .op(n11683) );
  nand4_1 U11283 ( .ip1(n11563), .ip2(n11562), .ip3(n11561), .ip4(n11560), 
        .op(n11564) );
  nor4_1 U11284 ( .ip1(n11593), .ip2(n11592), .ip3(n11591), .ip4(n11590), .op(
        n11594) );
  nand4_1 U11285 ( .ip1(n11585), .ip2(n11584), .ip3(n11583), .ip4(n11582), 
        .op(n11591) );
  nand4_1 U11286 ( .ip1(n11589), .ip2(n11588), .ip3(n11587), .ip4(n11586), 
        .op(n11590) );
  nand4_1 U11287 ( .ip1(n11581), .ip2(n11580), .ip3(n11579), .ip4(n11578), 
        .op(n11592) );
  and2_1 U11288 ( .ip1(n11955), .ip2(n11954), .op(n13575) );
  nand2_1 U11289 ( .ip1(n11927), .ip2(n13570), .op(n11955) );
  nand3_1 U11290 ( .ip1(n13741), .ip2(n13740), .ip3(n13739), .op(n13749) );
  nor2_1 U11291 ( .ip1(n13611), .ip2(n10223), .op(n13612) );
  inv_1 U11292 ( .ip(n16525), .op(n13611) );
  nand2_1 U11293 ( .ip1(n10194), .ip2(n10187), .op(n13911) );
  inv_1 U11294 ( .ip(n12932), .op(n17042) );
  and2_1 U11295 ( .ip1(n10193), .ip2(n17006), .op(n17007) );
  nand4_1 U11296 ( .ip1(n16687), .ip2(n16686), .ip3(n16685), .ip4(n17524), 
        .op(n19439) );
  inv_1 U11297 ( .ip(n16494), .op(n16495) );
  nand4_1 U11298 ( .ip1(n16643), .ip2(n17488), .ip3(n16642), .ip4(n16641), 
        .op(n17542) );
  nand2_1 U11299 ( .ip1(n13853), .ip2(n13997), .op(n16900) );
  inv_1 U11300 ( .ip(n13908), .op(n13853) );
  inv_1 U11301 ( .ip(n13678), .op(n20221) );
  nand4_1 U11302 ( .ip1(n16850), .ip2(n16849), .ip3(n16848), .ip4(n16847), 
        .op(n17166) );
  nor4_1 U11303 ( .ip1(n17274), .ip2(n17273), .ip3(n17272), .ip4(n17271), .op(
        n19059) );
  nand2_1 U11304 ( .ip1(n13984), .ip2(n13779), .op(n19073) );
  inv_1 U11305 ( .ip(n19069), .op(n19067) );
  nand2_1 U11306 ( .ip1(n13975), .ip2(n13977), .op(n18924) );
  nand4_1 U11307 ( .ip1(n16942), .ip2(n16941), .ip3(n16940), .ip4(n16939), 
        .op(n17167) );
  inv_1 U11308 ( .ip(n10181), .op(n17073) );
  nor4_1 U11309 ( .ip1(n16589), .ip2(n16588), .ip3(n17486), .ip4(n16763), .op(
        n19422) );
  nand4_1 U11310 ( .ip1(n13459), .ip2(n13458), .ip3(n13457), .ip4(n13456), 
        .op(n13460) );
  nor4_1 U11311 ( .ip1(n13514), .ip2(n13513), .ip3(n13512), .ip4(n13511), .op(
        n13515) );
  nand4_1 U11312 ( .ip1(n13502), .ip2(n13501), .ip3(n13500), .ip4(n13499), 
        .op(n13512) );
  nand4_1 U11313 ( .ip1(n13510), .ip2(n13509), .ip3(n13508), .ip4(n13507), 
        .op(n13511) );
  nand4_1 U11314 ( .ip1(n13494), .ip2(n13493), .ip3(n13492), .ip4(n13491), 
        .op(n13513) );
  nand2_1 U11315 ( .ip1(n14166), .ip2(n14165), .op(n14168) );
  and2_1 U11316 ( .ip1(n14169), .ip2(n17888), .op(n14241) );
  nand2_1 U11317 ( .ip1(n14213), .ip2(n14212), .op(n17987) );
  nor2_1 U11318 ( .ip1(n21161), .ip2(n14196), .op(n14197) );
  nand2_1 U11319 ( .ip1(n14262), .ip2(n14291), .op(n14579) );
  xnor2_1 U11320 ( .ip1(n14351), .ip2(n14350), .op(n14358) );
  nand2_2 U11321 ( .ip1(n14241), .ip2(n10372), .op(n14392) );
  nor2_1 U11322 ( .ip1(n14481), .ip2(n14434), .op(n14482) );
  nor2_1 U11323 ( .ip1(n14546), .ip2(n14485), .op(n14481) );
  nand4_1 U11324 ( .ip1(n12055), .ip2(n12054), .ip3(n12053), .ip4(n12052), 
        .op(n12056) );
  nor4_1 U11325 ( .ip1(n12085), .ip2(n12084), .ip3(n12083), .ip4(n12082), .op(
        n12086) );
  nand4_1 U11326 ( .ip1(n12077), .ip2(n12076), .ip3(n12075), .ip4(n12074), 
        .op(n12083) );
  nand4_1 U11327 ( .ip1(n12069), .ip2(n12068), .ip3(n12067), .ip4(n12066), 
        .op(n12085) );
  nand4_1 U11328 ( .ip1(n12081), .ip2(n12080), .ip3(n12079), .ip4(n12078), 
        .op(n12082) );
  nand4_1 U11329 ( .ip1(n10662), .ip2(n10661), .ip3(n10660), .ip4(n10659), 
        .op(n10663) );
  nor4_1 U11330 ( .ip1(n10692), .ip2(n10691), .ip3(n10690), .ip4(n10689), .op(
        n10693) );
  nand4_1 U11331 ( .ip1(n10684), .ip2(n10683), .ip3(n10682), .ip4(n10681), 
        .op(n10690) );
  nand4_1 U11332 ( .ip1(n10676), .ip2(n10675), .ip3(n10674), .ip4(n10673), 
        .op(n10692) );
  nand4_1 U11333 ( .ip1(n10688), .ip2(n10687), .ip3(n10686), .ip4(n10685), 
        .op(n10689) );
  nand4_1 U11334 ( .ip1(n12193), .ip2(n12192), .ip3(n12191), .ip4(n12190), 
        .op(n12194) );
  nor4_1 U11335 ( .ip1(n12223), .ip2(n12222), .ip3(n12221), .ip4(n12220), .op(
        n12224) );
  nand4_1 U11336 ( .ip1(n12215), .ip2(n12214), .ip3(n12213), .ip4(n12212), 
        .op(n12221) );
  nand4_1 U11337 ( .ip1(n12207), .ip2(n12206), .ip3(n12205), .ip4(n12204), 
        .op(n12223) );
  nand4_1 U11338 ( .ip1(n12219), .ip2(n12218), .ip3(n12217), .ip4(n12216), 
        .op(n12220) );
  nand4_1 U11339 ( .ip1(n12283), .ip2(n12282), .ip3(n12281), .ip4(n12280), 
        .op(n12284) );
  nor4_1 U11340 ( .ip1(n12313), .ip2(n12312), .ip3(n12311), .ip4(n12310), .op(
        n12314) );
  nand4_1 U11341 ( .ip1(n12305), .ip2(n12304), .ip3(n12303), .ip4(n12302), 
        .op(n12311) );
  nand4_1 U11342 ( .ip1(n12297), .ip2(n12296), .ip3(n12295), .ip4(n12294), 
        .op(n12313) );
  nand4_1 U11343 ( .ip1(n12309), .ip2(n12308), .ip3(n12307), .ip4(n12306), 
        .op(n12310) );
  nand4_1 U11344 ( .ip1(n11331), .ip2(n11330), .ip3(n11329), .ip4(n11328), 
        .op(n11332) );
  nor4_1 U11345 ( .ip1(n11361), .ip2(n11360), .ip3(n11359), .ip4(n11358), .op(
        n11362) );
  nand4_1 U11346 ( .ip1(n11353), .ip2(n11352), .ip3(n11351), .ip4(n11350), 
        .op(n11359) );
  nand4_1 U11347 ( .ip1(n11345), .ip2(n11344), .ip3(n11343), .ip4(n11342), 
        .op(n11361) );
  nand4_1 U11348 ( .ip1(n11357), .ip2(n11356), .ip3(n11355), .ip4(n11354), 
        .op(n11358) );
  nand4_1 U11349 ( .ip1(n11790), .ip2(n11789), .ip3(n11788), .ip4(n11787), 
        .op(n11791) );
  nor4_1 U11350 ( .ip1(n11820), .ip2(n11819), .ip3(n11818), .ip4(n11817), .op(
        n11821) );
  nand4_1 U11351 ( .ip1(n11812), .ip2(n11811), .ip3(n11810), .ip4(n11809), 
        .op(n11818) );
  nand4_1 U11352 ( .ip1(n11804), .ip2(n11803), .ip3(n11802), .ip4(n11801), 
        .op(n11820) );
  nand4_1 U11353 ( .ip1(n11816), .ip2(n11815), .ip3(n11814), .ip4(n11813), 
        .op(n11817) );
  inv_1 U11354 ( .ip(n18040), .op(n11784) );
  nand4_1 U11355 ( .ip1(n11606), .ip2(n11605), .ip3(n11604), .ip4(n11603), 
        .op(n11607) );
  nor4_1 U11356 ( .ip1(n11636), .ip2(n11635), .ip3(n11634), .ip4(n11633), .op(
        n11637) );
  nand4_1 U11357 ( .ip1(n11628), .ip2(n11627), .ip3(n11626), .ip4(n11625), 
        .op(n11634) );
  nand4_1 U11358 ( .ip1(n11620), .ip2(n11619), .ip3(n11618), .ip4(n11617), 
        .op(n11636) );
  nand4_1 U11359 ( .ip1(n11632), .ip2(n11631), .ip3(n11630), .ip4(n11629), 
        .op(n11633) );
  nand4_1 U11360 ( .ip1(n10354), .ip2(n14596), .ip3(n10353), .ip4(n22120), 
        .op(n10355) );
  nand4_1 U11361 ( .ip1(n13161), .ip2(n13160), .ip3(n13159), .ip4(n13158), 
        .op(n13163) );
  nand4_1 U11362 ( .ip1(n12928), .ip2(n12927), .ip3(n12926), .ip4(n12925), 
        .op(n12929) );
  nand4_1 U11363 ( .ip1(n13381), .ip2(n13380), .ip3(n13379), .ip4(n13378), 
        .op(n13382) );
  nor4_1 U11364 ( .ip1(n13436), .ip2(n13435), .ip3(n13434), .ip4(n13433), .op(
        n13437) );
  nand4_1 U11365 ( .ip1(n13424), .ip2(n13423), .ip3(n13422), .ip4(n13421), 
        .op(n13434) );
  nand4_1 U11366 ( .ip1(n13408), .ip2(n13407), .ip3(n13406), .ip4(n13405), 
        .op(n13436) );
  nand4_1 U11367 ( .ip1(n13432), .ip2(n13431), .ip3(n13430), .ip4(n13429), 
        .op(n13433) );
  nand4_1 U11368 ( .ip1(n13280), .ip2(n13279), .ip3(n13278), .ip4(n13277), 
        .op(n13281) );
  nor4_1 U11369 ( .ip1(n13310), .ip2(n13309), .ip3(n13308), .ip4(n13307), .op(
        n13311) );
  nand4_1 U11370 ( .ip1(n13302), .ip2(n13301), .ip3(n13300), .ip4(n13299), 
        .op(n13308) );
  nand4_1 U11371 ( .ip1(n13294), .ip2(n13293), .ip3(n13292), .ip4(n13291), 
        .op(n13310) );
  nand4_1 U11372 ( .ip1(n13306), .ip2(n13305), .ip3(n13304), .ip4(n13303), 
        .op(n13307) );
  nor4_1 U11373 ( .ip1(n13206), .ip2(n13205), .ip3(n13204), .ip4(n13203), .op(
        n15290) );
  nand4_1 U11374 ( .ip1(n13182), .ip2(n13181), .ip3(n13180), .ip4(n13179), 
        .op(n13204) );
  nand4_1 U11375 ( .ip1(n13178), .ip2(n13177), .ip3(n13176), .ip4(n13175), 
        .op(n13205) );
  nand4_1 U11376 ( .ip1(n13078), .ip2(n13077), .ip3(n13076), .ip4(n13075), 
        .op(n13079) );
  nor4_1 U11377 ( .ip1(n13108), .ip2(n13107), .ip3(n13106), .ip4(n13105), .op(
        n13109) );
  nand4_1 U11378 ( .ip1(n13100), .ip2(n13099), .ip3(n13098), .ip4(n13097), 
        .op(n13106) );
  nand4_1 U11379 ( .ip1(n13092), .ip2(n13091), .ip3(n13090), .ip4(n13089), 
        .op(n13108) );
  nand4_1 U11380 ( .ip1(n13104), .ip2(n13103), .ip3(n13102), .ip4(n13101), 
        .op(n13105) );
  inv_1 U11381 ( .ip(n17900), .op(n13072) );
  nand2_1 U11382 ( .ip1(n12880), .ip2(n17931), .op(n17296) );
  nand4_1 U11383 ( .ip1(n12879), .ip2(n12878), .ip3(n12877), .ip4(n12876), 
        .op(n12881) );
  nand4_1 U11384 ( .ip1(n12748), .ip2(n12747), .ip3(n12746), .ip4(n12745), 
        .op(n12749) );
  nor4_1 U11385 ( .ip1(n12778), .ip2(n12777), .ip3(n12776), .ip4(n12775), .op(
        n12779) );
  nand4_1 U11386 ( .ip1(n12770), .ip2(n12769), .ip3(n12768), .ip4(n12767), 
        .op(n12776) );
  nand4_1 U11387 ( .ip1(n12762), .ip2(n12761), .ip3(n12760), .ip4(n12759), 
        .op(n12778) );
  nand4_1 U11388 ( .ip1(n12774), .ip2(n12773), .ip3(n12772), .ip4(n12771), 
        .op(n12775) );
  nand4_1 U11389 ( .ip1(n12938), .ip2(n12937), .ip3(n12936), .ip4(n12935), 
        .op(n12939) );
  nor4_1 U11390 ( .ip1(n12968), .ip2(n12967), .ip3(n12966), .ip4(n12965), .op(
        n12969) );
  nand4_1 U11391 ( .ip1(n12960), .ip2(n12959), .ip3(n12958), .ip4(n12957), 
        .op(n12966) );
  nand4_1 U11392 ( .ip1(n12952), .ip2(n12951), .ip3(n12950), .ip4(n12949), 
        .op(n12968) );
  nand4_1 U11393 ( .ip1(n12964), .ip2(n12963), .ip3(n12962), .ip4(n12961), 
        .op(n12965) );
  nand4_1 U11394 ( .ip1(n13018), .ip2(n13017), .ip3(n13016), .ip4(n13015), 
        .op(n13019) );
  nand4_1 U11395 ( .ip1(n13028), .ip2(n13027), .ip3(n13026), .ip4(n13025), 
        .op(n13029) );
  nor4_1 U11396 ( .ip1(n13058), .ip2(n13057), .ip3(n13056), .ip4(n13055), .op(
        n13059) );
  nand4_1 U11397 ( .ip1(n13050), .ip2(n13049), .ip3(n13048), .ip4(n13047), 
        .op(n13056) );
  nand4_1 U11398 ( .ip1(n13042), .ip2(n13041), .ip3(n13040), .ip4(n13039), 
        .op(n13058) );
  nand4_1 U11399 ( .ip1(n13054), .ip2(n13053), .ip3(n13052), .ip4(n13051), 
        .op(n13055) );
  nand4_1 U11400 ( .ip1(n12639), .ip2(n12638), .ip3(n12637), .ip4(n12636), 
        .op(n12640) );
  nand4_1 U11401 ( .ip1(n12557), .ip2(n12556), .ip3(n12555), .ip4(n12554), 
        .op(n12558) );
  nor4_1 U11402 ( .ip1(n12587), .ip2(n12586), .ip3(n12585), .ip4(n12584), .op(
        n12588) );
  nand4_1 U11403 ( .ip1(n12579), .ip2(n12578), .ip3(n12577), .ip4(n12576), 
        .op(n12585) );
  nand4_1 U11404 ( .ip1(n12571), .ip2(n12570), .ip3(n12569), .ip4(n12568), 
        .op(n12587) );
  nand4_1 U11405 ( .ip1(n12583), .ip2(n12582), .ip3(n12581), .ip4(n12580), 
        .op(n12584) );
  nand4_1 U11406 ( .ip1(n12648), .ip2(n12647), .ip3(n12646), .ip4(n12645), 
        .op(n12649) );
  nor4_1 U11407 ( .ip1(n12678), .ip2(n12677), .ip3(n12676), .ip4(n12675), .op(
        n12679) );
  nand4_1 U11408 ( .ip1(n12670), .ip2(n12669), .ip3(n12668), .ip4(n12667), 
        .op(n12676) );
  nand4_1 U11409 ( .ip1(n12662), .ip2(n12661), .ip3(n12660), .ip4(n12659), 
        .op(n12678) );
  nand4_1 U11410 ( .ip1(n12674), .ip2(n12673), .ip3(n12672), .ip4(n12671), 
        .op(n12675) );
  nand4_1 U11411 ( .ip1(n12702), .ip2(n12701), .ip3(n12700), .ip4(n12699), 
        .op(n12703) );
  nor4_1 U11412 ( .ip1(n12732), .ip2(n12731), .ip3(n12730), .ip4(n12729), .op(
        n12733) );
  nand4_1 U11413 ( .ip1(n12724), .ip2(n12723), .ip3(n12722), .ip4(n12721), 
        .op(n12730) );
  nand4_1 U11414 ( .ip1(n12728), .ip2(n12727), .ip3(n12726), .ip4(n12725), 
        .op(n12729) );
  nand4_1 U11415 ( .ip1(n12720), .ip2(n12719), .ip3(n12718), .ip4(n12717), 
        .op(n12731) );
  nand4_1 U11416 ( .ip1(n13363), .ip2(n13362), .ip3(n13361), .ip4(n13360), 
        .op(n13365) );
  nand2_1 U11417 ( .ip1(n13266), .ip2(n13265), .op(n15789) );
  nand2_1 U11418 ( .ip1(n13264), .ip2(n10200), .op(n13266) );
  or2_1 U11419 ( .ip1(n10200), .ip2(n15291), .op(n13265) );
  nand4_1 U11420 ( .ip1(n13263), .ip2(n13262), .ip3(n13261), .ip4(n13260), 
        .op(n13264) );
  nand4_1 U11421 ( .ip1(n12378), .ip2(n12377), .ip3(n12376), .ip4(n12375), 
        .op(n12379) );
  nor4_1 U11422 ( .ip1(n12408), .ip2(n12407), .ip3(n12406), .ip4(n12405), .op(
        n12409) );
  nand4_1 U11423 ( .ip1(n12400), .ip2(n12399), .ip3(n12398), .ip4(n12397), 
        .op(n12406) );
  nand4_1 U11424 ( .ip1(n12392), .ip2(n12391), .ip3(n12390), .ip4(n12389), 
        .op(n12408) );
  nand4_1 U11425 ( .ip1(n12404), .ip2(n12403), .ip3(n12402), .ip4(n12401), 
        .op(n12405) );
  nand4_1 U11426 ( .ip1(n12467), .ip2(n12466), .ip3(n12465), .ip4(n12464), 
        .op(n12468) );
  nor4_1 U11427 ( .ip1(n12497), .ip2(n12496), .ip3(n12495), .ip4(n12494), .op(
        n12498) );
  nand4_1 U11428 ( .ip1(n12489), .ip2(n12488), .ip3(n12487), .ip4(n12486), 
        .op(n12495) );
  nand4_1 U11429 ( .ip1(n12481), .ip2(n12480), .ip3(n12479), .ip4(n12478), 
        .op(n12497) );
  nand4_1 U11430 ( .ip1(n12493), .ip2(n12492), .ip3(n12491), .ip4(n12490), 
        .op(n12494) );
  nand4_1 U11431 ( .ip1(n12008), .ip2(n12007), .ip3(n12006), .ip4(n12005), 
        .op(n12009) );
  nor4_1 U11432 ( .ip1(n12038), .ip2(n12037), .ip3(n12036), .ip4(n12035), .op(
        n12039) );
  nand4_1 U11433 ( .ip1(n12030), .ip2(n12029), .ip3(n12028), .ip4(n12027), 
        .op(n12036) );
  nand4_1 U11434 ( .ip1(n12022), .ip2(n12021), .ip3(n12020), .ip4(n12019), 
        .op(n12038) );
  nand4_1 U11435 ( .ip1(n12034), .ip2(n12033), .ip3(n12032), .ip4(n12031), 
        .op(n12035) );
  nand4_1 U11436 ( .ip1(n12134), .ip2(n12133), .ip3(n12132), .ip4(n12131), 
        .op(n12135) );
  nand4_1 U11437 ( .ip1(n12831), .ip2(n12830), .ip3(n12829), .ip4(n12828), 
        .op(n12832) );
  nand4_1 U11438 ( .ip1(n10433), .ip2(n10432), .ip3(n10431), .ip4(n10430), 
        .op(n10445) );
  nand4_1 U11439 ( .ip1(n10753), .ip2(n10752), .ip3(n10751), .ip4(n10750), 
        .op(n10754) );
  nor4_1 U11440 ( .ip1(n10783), .ip2(n10782), .ip3(n10781), .ip4(n10780), .op(
        n10784) );
  nand4_1 U11441 ( .ip1(n10775), .ip2(n10774), .ip3(n10773), .ip4(n10772), 
        .op(n10781) );
  nand4_1 U11442 ( .ip1(n10767), .ip2(n10766), .ip3(n10765), .ip4(n10764), 
        .op(n10783) );
  nand4_1 U11443 ( .ip1(n10779), .ip2(n10778), .ip3(n10777), .ip4(n10776), 
        .op(n10780) );
  nand4_1 U11444 ( .ip1(n10569), .ip2(n10568), .ip3(n10567), .ip4(n10566), 
        .op(n10570) );
  nor4_1 U11445 ( .ip1(n10599), .ip2(n10598), .ip3(n10597), .ip4(n10596), .op(
        n10600) );
  nand4_1 U11446 ( .ip1(n10591), .ip2(n10590), .ip3(n10589), .ip4(n10588), 
        .op(n10597) );
  nand4_1 U11447 ( .ip1(n10583), .ip2(n10582), .ip3(n10581), .ip4(n10580), 
        .op(n10599) );
  nand4_1 U11448 ( .ip1(n10595), .ip2(n10594), .ip3(n10593), .ip4(n10592), 
        .op(n10596) );
  nand4_1 U11449 ( .ip1(n10461), .ip2(n10460), .ip3(n10459), .ip4(n10458), 
        .op(n10462) );
  nor4_1 U11450 ( .ip1(n10503), .ip2(n10502), .ip3(n10501), .ip4(n10500), .op(
        n10504) );
  nand4_1 U11451 ( .ip1(n10491), .ip2(n10490), .ip3(n10489), .ip4(n10488), 
        .op(n10501) );
  nand4_1 U11452 ( .ip1(n10479), .ip2(n10478), .ip3(n10477), .ip4(n10476), 
        .op(n10503) );
  nand4_1 U11453 ( .ip1(n10499), .ip2(n10498), .ip3(n10497), .ip4(n10496), 
        .op(n10500) );
  inv_1 U11454 ( .ip(n18579), .op(n10455) );
  nand4_1 U11455 ( .ip1(n10526), .ip2(n10525), .ip3(n10524), .ip4(n10523), 
        .op(n10527) );
  nor4_1 U11456 ( .ip1(n10556), .ip2(n10555), .ip3(n10554), .ip4(n10553), .op(
        n10557) );
  nand4_1 U11457 ( .ip1(n10548), .ip2(n10547), .ip3(n10546), .ip4(n10545), 
        .op(n10554) );
  nand4_1 U11458 ( .ip1(n10552), .ip2(n10551), .ip3(n10550), .ip4(n10549), 
        .op(n10553) );
  nand4_1 U11459 ( .ip1(n10544), .ip2(n10543), .ip3(n10542), .ip4(n10541), 
        .op(n10555) );
  nand4_1 U11460 ( .ip1(n11413), .ip2(n11412), .ip3(n11411), .ip4(n11410), 
        .op(n11414) );
  nand4_1 U11461 ( .ip1(n11043), .ip2(n11042), .ip3(n11041), .ip4(n11040), 
        .op(n11044) );
  nor4_1 U11462 ( .ip1(n11073), .ip2(n11072), .ip3(n11071), .ip4(n11070), .op(
        n11074) );
  nand4_1 U11463 ( .ip1(n11065), .ip2(n11064), .ip3(n11063), .ip4(n11062), 
        .op(n11071) );
  nand4_1 U11464 ( .ip1(n11057), .ip2(n11056), .ip3(n11055), .ip4(n11054), 
        .op(n11073) );
  nand4_1 U11465 ( .ip1(n11069), .ip2(n11068), .ip3(n11067), .ip4(n11066), 
        .op(n11070) );
  nand4_1 U11466 ( .ip1(n10891), .ip2(n10890), .ip3(n10889), .ip4(n10888), 
        .op(n17398) );
  nor4_1 U11467 ( .ip1(n10887), .ip2(n10886), .ip3(n10885), .ip4(n10884), .op(
        n10888) );
  nand2_1 U11468 ( .ip1(n10985), .ip2(n17399), .op(n17404) );
  nand4_1 U11469 ( .ip1(n11514), .ip2(n11513), .ip3(n11512), .ip4(n11511), 
        .op(n11515) );
  nor4_1 U11470 ( .ip1(n11544), .ip2(n11543), .ip3(n11542), .ip4(n11541), .op(
        n11545) );
  nand4_1 U11471 ( .ip1(n11536), .ip2(n11535), .ip3(n11534), .ip4(n11533), 
        .op(n11542) );
  nand4_1 U11472 ( .ip1(n11528), .ip2(n11527), .ip3(n11526), .ip4(n11525), 
        .op(n11544) );
  nand4_1 U11473 ( .ip1(n11540), .ip2(n11539), .ip3(n11538), .ip4(n11537), 
        .op(n11541) );
  mux2_2 U11474 ( .ip1(n18341), .ip2(n11457), .s(n12683), .op(n21282) );
  nand4_1 U11475 ( .ip1(n11456), .ip2(n11455), .ip3(n11454), .ip4(n11453), 
        .op(n11457) );
  nand4_1 U11476 ( .ip1(n10619), .ip2(n10618), .ip3(n10617), .ip4(n10616), 
        .op(n10620) );
  nor4_1 U11477 ( .ip1(n10649), .ip2(n10648), .ip3(n10647), .ip4(n10646), .op(
        n10650) );
  nand4_1 U11478 ( .ip1(n10641), .ip2(n10640), .ip3(n10639), .ip4(n10638), 
        .op(n10647) );
  nand4_1 U11479 ( .ip1(n10645), .ip2(n10644), .ip3(n10643), .ip4(n10642), 
        .op(n10646) );
  nand4_1 U11480 ( .ip1(n10637), .ip2(n10636), .ip3(n10635), .ip4(n10634), 
        .op(n10648) );
  nand4_1 U11481 ( .ip1(n12149), .ip2(n12148), .ip3(n12147), .ip4(n12146), 
        .op(n12150) );
  nor4_1 U11482 ( .ip1(n12179), .ip2(n12178), .ip3(n12177), .ip4(n12176), .op(
        n12180) );
  nand4_1 U11483 ( .ip1(n12171), .ip2(n12170), .ip3(n12169), .ip4(n12168), 
        .op(n12177) );
  nand4_1 U11484 ( .ip1(n12175), .ip2(n12174), .ip3(n12173), .ip4(n12172), 
        .op(n12176) );
  nand4_1 U11485 ( .ip1(n12167), .ip2(n12166), .ip3(n12165), .ip4(n12164), 
        .op(n12178) );
  nand4_1 U11486 ( .ip1(n12274), .ip2(n12273), .ip3(n12272), .ip4(n12271), 
        .op(n12275) );
  nand4_1 U11487 ( .ip1(n11125), .ip2(n11124), .ip3(n11123), .ip4(n11122), 
        .op(n11126) );
  nand4_1 U11488 ( .ip1(n11031), .ip2(n11030), .ip3(n11029), .ip4(n11028), 
        .op(n11035) );
  nand4_1 U11489 ( .ip1(n11288), .ip2(n11287), .ip3(n11286), .ip4(n11285), 
        .op(n11289) );
  nor4_1 U11490 ( .ip1(n11318), .ip2(n11317), .ip3(n11316), .ip4(n11315), .op(
        n11319) );
  nand4_1 U11491 ( .ip1(n11310), .ip2(n11309), .ip3(n11308), .ip4(n11307), 
        .op(n11316) );
  nand4_1 U11492 ( .ip1(n11314), .ip2(n11313), .ip3(n11312), .ip4(n11311), 
        .op(n11315) );
  nand4_1 U11493 ( .ip1(n11306), .ip2(n11305), .ip3(n11304), .ip4(n11303), 
        .op(n11317) );
  nand4_1 U11494 ( .ip1(n11746), .ip2(n11745), .ip3(n11744), .ip4(n11743), 
        .op(n11747) );
  nor4_1 U11495 ( .ip1(n11776), .ip2(n11775), .ip3(n11774), .ip4(n11773), .op(
        n11777) );
  nand4_1 U11496 ( .ip1(n11768), .ip2(n11767), .ip3(n11766), .ip4(n11765), 
        .op(n11774) );
  nand4_1 U11497 ( .ip1(n11772), .ip2(n11771), .ip3(n11770), .ip4(n11769), 
        .op(n11773) );
  nand4_1 U11498 ( .ip1(n11764), .ip2(n11763), .ip3(n11762), .ip4(n11761), 
        .op(n11775) );
  nand4_1 U11499 ( .ip1(n11275), .ip2(n11274), .ip3(n11273), .ip4(n11272), 
        .op(n11276) );
  nand4_1 U11500 ( .ip1(n11917), .ip2(n11916), .ip3(n11915), .ip4(n11914), 
        .op(n11918) );
  nor4_1 U11501 ( .ip1(n11913), .ip2(n11912), .ip3(n11911), .ip4(n11910), .op(
        n11914) );
  nand4_1 U11502 ( .ip1(n11232), .ip2(n11231), .ip3(n11230), .ip4(n11229), 
        .op(n11233) );
  nand4_1 U11503 ( .ip1(n12458), .ip2(n12457), .ip3(n12456), .ip4(n12455), 
        .op(n12459) );
  nand4_1 U11504 ( .ip1(n12369), .ip2(n12368), .ip3(n12367), .ip4(n12366), 
        .op(n12370) );
  nand4_1 U11505 ( .ip1(n11873), .ip2(n11872), .ip3(n11871), .ip4(n11870), 
        .op(n11874) );
  nand4_1 U11506 ( .ip1(n11470), .ip2(n11469), .ip3(n11468), .ip4(n11467), 
        .op(n11471) );
  nor4_1 U11507 ( .ip1(n11500), .ip2(n11499), .ip3(n11498), .ip4(n11497), .op(
        n11501) );
  nand4_1 U11508 ( .ip1(n11492), .ip2(n11491), .ip3(n11490), .ip4(n11489), 
        .op(n11498) );
  nand4_1 U11509 ( .ip1(n11496), .ip2(n11495), .ip3(n11494), .ip4(n11493), 
        .op(n11497) );
  nand4_1 U11510 ( .ip1(n11488), .ip2(n11487), .ip3(n11486), .ip4(n11485), 
        .op(n11499) );
  nand4_1 U11511 ( .ip1(n11998), .ip2(n11997), .ip3(n11996), .ip4(n11995), 
        .op(n12000) );
  nand4_1 U11512 ( .ip1(n10743), .ip2(n10742), .ip3(n10741), .ip4(n10740), 
        .op(n10744) );
  nand4_1 U11513 ( .ip1(n15330), .ip2(n10354), .ip3(n22112), .ip4(n15339), 
        .op(n10343) );
  nand4_1 U11514 ( .ip1(n11697), .ip2(n11696), .ip3(n11695), .ip4(n11694), 
        .op(n11698) );
  nor4_1 U11515 ( .ip1(n11727), .ip2(n11726), .ip3(n11725), .ip4(n11724), .op(
        n11728) );
  nand4_1 U11516 ( .ip1(n11719), .ip2(n11718), .ip3(n11717), .ip4(n11716), 
        .op(n11725) );
  nand4_1 U11517 ( .ip1(n11711), .ip2(n11710), .ip3(n11709), .ip4(n11708), 
        .op(n11727) );
  nand4_1 U11518 ( .ip1(n11723), .ip2(n11722), .ip3(n11721), .ip4(n11720), 
        .op(n11724) );
  inv_1 U11519 ( .ip(n21584), .op(n11691) );
  nand4_1 U11520 ( .ip1(n11653), .ip2(n11652), .ip3(n11651), .ip4(n11650), 
        .op(n11654) );
  nor4_1 U11521 ( .ip1(n11683), .ip2(n11682), .ip3(n11681), .ip4(n11680), .op(
        n11684) );
  nand4_1 U11522 ( .ip1(n11675), .ip2(n11674), .ip3(n11673), .ip4(n11672), 
        .op(n11681) );
  nand4_1 U11523 ( .ip1(n11679), .ip2(n11678), .ip3(n11677), .ip4(n11676), 
        .op(n11680) );
  nand4_1 U11524 ( .ip1(n11671), .ip2(n11670), .ip3(n11669), .ip4(n11668), 
        .op(n11682) );
  nand4_1 U11525 ( .ip1(n11597), .ip2(n11596), .ip3(n11595), .ip4(n11594), 
        .op(n11598) );
  nand4_1 U11526 ( .ip1(n21539), .ip2(n19427), .ip3(n21538), .ip4(n21537), 
        .op(n21543) );
  nand4_1 U11527 ( .ip1(n20235), .ip2(n20234), .ip3(n20233), .ip4(n20232), 
        .op(n20236) );
  nand4_1 U11528 ( .ip1(n17538), .ip2(n17537), .ip3(n17536), .ip4(n17535), 
        .op(n17539) );
  nand4_1 U11529 ( .ip1(n18377), .ip2(n18748), .ip3(n18376), .ip4(n18375), 
        .op(n18380) );
  nor4_1 U11530 ( .ip1(n18941), .ip2(n18940), .ip3(n18939), .ip4(n18938), .op(
        n18942) );
  nand4_1 U11531 ( .ip1(n13518), .ip2(n13517), .ip3(n13516), .ip4(n13515), 
        .op(n13519) );
  nor2_1 U11532 ( .ip1(n14292), .ip2(n14291), .op(n20692) );
  nand2_1 U11533 ( .ip1(n14363), .ip2(n14364), .op(n17431) );
  nand2_1 U11534 ( .ip1(n14298), .ip2(n14586), .op(n14307) );
  nand2_1 U11535 ( .ip1(n14355), .ip2(n14354), .op(n18294) );
  nor2_1 U11536 ( .ip1(n14357), .ip2(n14358), .op(n20021) );
  nand2_1 U11537 ( .ip1(n14512), .ip2(n14511), .op(n14513) );
  and2_1 U11538 ( .ip1(n14047), .ip2(n14046), .op(n14503) );
  nand2_1 U11539 ( .ip1(n14536), .ip2(n14535), .op(n14544) );
  inv_1 U11540 ( .ip(n14573), .op(n14536) );
  inv_1 U11541 ( .ip(n14560), .op(n14557) );
  nand2_1 U11542 ( .ip1(n14550), .ip2(n14549), .op(n14554) );
  nand2_1 U11543 ( .ip1(n14536), .ip2(n14552), .op(n14553) );
  nor2_1 U11544 ( .ip1(n14562), .ip2(n14561), .op(n14563) );
  inv_1 U11545 ( .ip(n14558), .op(n14562) );
  nor2_1 U11546 ( .ip1(n14560), .ip2(n10208), .op(n14561) );
  mux2_2 U11547 ( .ip1(n19330), .ip2(n12090), .s(n13315), .op(n22064) );
  nand4_1 U11548 ( .ip1(n12089), .ip2(n12088), .ip3(n12087), .ip4(n12086), 
        .op(n12090) );
  nand4_1 U11549 ( .ip1(n10696), .ip2(n10695), .ip3(n10694), .ip4(n10693), 
        .op(n10697) );
  mux2_2 U11550 ( .ip1(n19342), .ip2(n12228), .s(n13315), .op(n22062) );
  nand4_1 U11551 ( .ip1(n12227), .ip2(n12226), .ip3(n12225), .ip4(n12224), 
        .op(n12228) );
  nand4_1 U11552 ( .ip1(n12317), .ip2(n12316), .ip3(n12315), .ip4(n12314), 
        .op(n12318) );
  mux2_2 U11553 ( .ip1(n19089), .ip2(n11366), .s(n13315), .op(n21281) );
  nand4_1 U11554 ( .ip1(n11365), .ip2(n11364), .ip3(n11363), .ip4(n11362), 
        .op(n11366) );
  nand2_1 U11555 ( .ip1(n11827), .ip2(n11826), .op(n22063) );
  nand4_1 U11556 ( .ip1(n11824), .ip2(n11823), .ip3(n11822), .ip4(n11821), 
        .op(n11825) );
  mux2_2 U11557 ( .ip1(n18867), .ip2(n11641), .s(n13315), .op(n22066) );
  nand4_1 U11558 ( .ip1(n11640), .ip2(n11639), .ip3(n11638), .ip4(n11637), 
        .op(n11641) );
  nand4_1 U11559 ( .ip1(n13440), .ip2(n13439), .ip3(n13438), .ip4(n13437), 
        .op(n13442) );
  nand4_1 U11560 ( .ip1(n13314), .ip2(n13313), .ip3(n13312), .ip4(n13311), 
        .op(n13316) );
  nand2_1 U11561 ( .ip1(n13113), .ip2(n13441), .op(n13114) );
  or2_1 U11562 ( .ip1(n13441), .ip2(n13072), .op(n13115) );
  nand4_1 U11563 ( .ip1(n13112), .ip2(n13111), .ip3(n13110), .ip4(n13109), 
        .op(n13113) );
  nand2_1 U11564 ( .ip1(n17297), .ip2(n17296), .op(n22061) );
  nand4_1 U11565 ( .ip1(n12782), .ip2(n12781), .ip3(n12780), .ip4(n12779), 
        .op(n12783) );
  mux2_2 U11566 ( .ip1(n18007), .ip2(n12973), .s(n13315), .op(n22065) );
  nand4_1 U11567 ( .ip1(n12972), .ip2(n12971), .ip3(n12970), .ip4(n12969), 
        .op(n12973) );
  nand4_1 U11568 ( .ip1(n13062), .ip2(n13061), .ip3(n13060), .ip4(n13059), 
        .op(n13064) );
  nand4_1 U11569 ( .ip1(n12591), .ip2(n12590), .ip3(n12589), .ip4(n12588), 
        .op(n12593) );
  mux2_1 U11570 ( .ip1(n18423), .ip2(n12684), .s(n12683), .op(n22054) );
  nand4_1 U11571 ( .ip1(n12682), .ip2(n12681), .ip3(n12680), .ip4(n12679), 
        .op(n12684) );
  nand4_1 U11572 ( .ip1(n12736), .ip2(n12735), .ip3(n12734), .ip4(n12733), 
        .op(n12737) );
  mux2_2 U11573 ( .ip1(n19396), .ip2(n12413), .s(n13315), .op(n22056) );
  nand4_1 U11574 ( .ip1(n12412), .ip2(n12411), .ip3(n12410), .ip4(n12409), 
        .op(n12413) );
  nand4_1 U11575 ( .ip1(n12501), .ip2(n12500), .ip3(n12499), .ip4(n12498), 
        .op(n12502) );
  mux2_2 U11576 ( .ip1(n18283), .ip2(n12043), .s(n13315), .op(n22068) );
  nand4_1 U11577 ( .ip1(n12042), .ip2(n12041), .ip3(n12040), .ip4(n12039), 
        .op(n12043) );
  nand4_1 U11578 ( .ip1(n10787), .ip2(n10786), .ip3(n10785), .ip4(n10784), 
        .op(n10788) );
  mux2_2 U11579 ( .ip1(n18515), .ip2(n10604), .s(n13315), .op(n22083) );
  nand4_1 U11580 ( .ip1(n10603), .ip2(n10602), .ip3(n10601), .ip4(n10600), 
        .op(n10604) );
  nand2_1 U11581 ( .ip1(n10510), .ip2(n10509), .op(n22084) );
  or2_1 U11582 ( .ip1(n12683), .ip2(n10455), .op(n10510) );
  nand4_1 U11583 ( .ip1(n10507), .ip2(n10506), .ip3(n10505), .ip4(n10504), 
        .op(n10508) );
  nand4_1 U11584 ( .ip1(n10560), .ip2(n10559), .ip3(n10558), .ip4(n10557), 
        .op(n10561) );
  nand4_1 U11585 ( .ip1(n11077), .ip2(n11076), .ip3(n11075), .ip4(n11074), 
        .op(n11078) );
  nand4_1 U11586 ( .ip1(n11548), .ip2(n11547), .ip3(n11546), .ip4(n11545), 
        .op(n11549) );
  nand4_1 U11587 ( .ip1(n10653), .ip2(n10652), .ip3(n10651), .ip4(n10650), 
        .op(n10654) );
  nand4_1 U11588 ( .ip1(n12183), .ip2(n12182), .ip3(n12181), .ip4(n12180), 
        .op(n12185) );
  nand4_1 U11589 ( .ip1(n11322), .ip2(n11321), .ip3(n11320), .ip4(n11319), 
        .op(n11323) );
  nand4_1 U11590 ( .ip1(n11780), .ip2(n11779), .ip3(n11778), .ip4(n11777), 
        .op(n11781) );
  nand2_1 U11591 ( .ip1(n11918), .ip2(n17399), .op(n11919) );
  inv_1 U11592 ( .ip(n19032), .op(n11877) );
  nand4_1 U11593 ( .ip1(n11504), .ip2(n11503), .ip3(n11502), .ip4(n11501), 
        .op(n11505) );
  nor4_1 U11594 ( .ip1(n15310), .ip2(n17883), .ip3(n10343), .ip4(n10342), .op(
        n17779) );
  nand2_1 U11595 ( .ip1(n11734), .ip2(n11733), .op(n22069) );
  or2_1 U11596 ( .ip1(n12683), .ip2(n11691), .op(n11734) );
  nand4_1 U11597 ( .ip1(n11731), .ip2(n11730), .ip3(n11729), .ip4(n11728), 
        .op(n11732) );
  nand4_1 U11598 ( .ip1(n11687), .ip2(n11686), .ip3(n11685), .ip4(n11684), 
        .op(n11688) );
  nand4_1 U11599 ( .ip1(n16749), .ip2(n16748), .ip3(n16747), .ip4(n16746), 
        .op(dmem_haddr[2]) );
  nand4_1 U11600 ( .ip1(n16787), .ip2(n16786), .ip3(n16785), .ip4(n16784), 
        .op(dmem_haddr[3]) );
  nand4_1 U11601 ( .ip1(n17242), .ip2(n17241), .ip3(n17240), .ip4(n17239), 
        .op(dmem_haddr[4]) );
  nand4_1 U11602 ( .ip1(n17072), .ip2(n17071), .ip3(n17070), .ip4(n17069), 
        .op(dmem_haddr[6]) );
  nand4_1 U11603 ( .ip1(n17019), .ip2(n17018), .ip3(n17017), .ip4(n17016), 
        .op(dmem_haddr[7]) );
  nand4_1 U11604 ( .ip1(n16823), .ip2(n16822), .ip3(n16821), .ip4(n16820), 
        .op(dmem_haddr[8]) );
  nand4_1 U11605 ( .ip1(n16986), .ip2(n16985), .ip3(n16984), .ip4(n16983), 
        .op(dmem_haddr[10]) );
  nand4_1 U11606 ( .ip1(n16703), .ip2(n16702), .ip3(n16701), .ip4(n16700), 
        .op(dmem_haddr[11]) );
  nand4_1 U11607 ( .ip1(n20741), .ip2(n20740), .ip3(n20739), .ip4(n20738), 
        .op(n20742) );
  nand4_1 U11608 ( .ip1(n17158), .ip2(n17157), .ip3(n17156), .ip4(n17155), 
        .op(dmem_haddr[14]) );
  nand4_1 U11609 ( .ip1(n16541), .ip2(n16540), .ip3(n16539), .ip4(n16538), 
        .op(dmem_haddr[16]) );
  nand4_1 U11610 ( .ip1(n16664), .ip2(n16663), .ip3(n16662), .ip4(n16661), 
        .op(dmem_haddr[17]) );
  nand4_1 U11611 ( .ip1(n16879), .ip2(n16878), .ip3(n16877), .ip4(n16876), 
        .op(dmem_haddr[18]) );
  nand4_1 U11612 ( .ip1(n16911), .ip2(n16910), .ip3(n16909), .ip4(n16908), 
        .op(dmem_haddr[19]) );
  nand4_1 U11613 ( .ip1(n17295), .ip2(n17294), .ip3(n17293), .ip4(n17292), 
        .op(dmem_haddr[20]) );
  nand4_1 U11614 ( .ip1(n17190), .ip2(n17189), .ip3(n17188), .ip4(n17187), 
        .op(dmem_haddr[22]) );
  nand4_1 U11615 ( .ip1(n16616), .ip2(n16615), .ip3(n16614), .ip4(n16613), 
        .op(dmem_haddr[23]) );
  nand4_1 U11616 ( .ip1(n16961), .ip2(n16960), .ip3(n16959), .ip4(n16958), 
        .op(dmem_haddr[26]) );
  nand4_1 U11617 ( .ip1(n17127), .ip2(n17126), .ip3(n17125), .ip4(n17124), 
        .op(dmem_haddr[30]) );
  nand2_1 U11618 ( .ip1(n14578), .ip2(n14302), .op(n20797) );
  inv_1 U11619 ( .ip(n14575), .op(n14576) );
  nand2_1 U11620 ( .ip1(n19893), .ip2(n14365), .op(n19896) );
  nand2_1 U11621 ( .ip1(n14523), .ip2(n14522), .op(n14524) );
  nand2_1 U11622 ( .ip1(n18285), .ip2(n18288), .op(n14523) );
  nand2_1 U11623 ( .ip1(n20038), .ip2(n19491), .op(n19492) );
  nand2_1 U11624 ( .ip1(n20042), .ip2(n20041), .op(n19491) );
  nand2_1 U11625 ( .ip1(n20044), .ip2(n20043), .op(n20045) );
  nor2_1 U11626 ( .ip1(n10183), .ip2(n20039), .op(n20044) );
  nand2_1 U11627 ( .ip1(n14573), .ip2(n14572), .op(n14574) );
  nand2_1 U11628 ( .ip1(n14528), .ip2(n14527), .op(n14529) );
  nand2_1 U11629 ( .ip1(n14475), .ip2(n14474), .op(n14492) );
  mux2_1 U11630 ( .ip1(dmem_hwdata[6]), .ip2(n22065), .s(n17777), .op(n8833)
         );
  mux2_1 U11631 ( .ip1(dmem_hwdata[7]), .ip2(n17376), .s(n17429), .op(n8832)
         );
  mux2_1 U11632 ( .ip1(\pipeline/store_data_WB [9]), .ip2(n22054), .s(n19498), 
        .op(n8830) );
  mux2_2 U11633 ( .ip1(dmem_hwdata[1]), .ip2(n22055), .s(n20389), .op(n8838)
         );
  mux2_1 U11634 ( .ip1(\pipeline/store_data_WB [15]), .ip2(n22068), .s(n22067), 
        .op(n8824) );
  mux2_1 U11635 ( .ip1(\pipeline/store_data_WB [14]), .ip2(n22064), .s(n22067), 
        .op(n8825) );
  mux2_1 U11636 ( .ip1(dmem_hwdata[4]), .ip2(n22061), .s(n17429), .op(n8835)
         );
  mux2_1 U11637 ( .ip1(\pipeline/store_data_WB [19]), .ip2(n22084), .s(n17429), 
        .op(n8820) );
  mux2_1 U11638 ( .ip1(\pipeline/store_data_WB [18]), .ip2(n22083), .s(n17777), 
        .op(n8821) );
  mux2_1 U11639 ( .ip1(\pipeline/store_data_WB [13]), .ip2(n22062), .s(n19498), 
        .op(n8826) );
  mux2_1 U11640 ( .ip1(\pipeline/store_data_WB [8]), .ip2(n22052), .s(n17777), 
        .op(n8831) );
  mux2_1 U11641 ( .ip1(\pipeline/store_data_WB [20]), .ip2(n22085), .s(n17777), 
        .op(n8819) );
  mux2_1 U11642 ( .ip1(\pipeline/store_data_WB [12]), .ip2(n22060), .s(n22067), 
        .op(n8827) );
  mux2_1 U11643 ( .ip1(\pipeline/store_data_WB [10]), .ip2(n22056), .s(n17777), 
        .op(n8829) );
  mux2_1 U11644 ( .ip1(\pipeline/store_data_WB [11]), .ip2(n22058), .s(n22067), 
        .op(n8828) );
  mux2_1 U11645 ( .ip1(\pipeline/store_data_WB [30]), .ip2(n22066), .s(n19498), 
        .op(n8809) );
  mux2_1 U11646 ( .ip1(\pipeline/store_data_WB [16]), .ip2(n22082), .s(n19498), 
        .op(n8823) );
  nand2_1 U11647 ( .ip1(imem_haddr[26]), .ip2(n21995), .op(n18346) );
  nand2_1 U11648 ( .ip1(n21995), .ip2(imem_haddr[23]), .op(n20107) );
  xor2_1 U11649 ( .ip1(n14493), .ip2(n14532), .op(imem_haddr[25]) );
  nand2_1 U11650 ( .ip1(n14563), .ip2(n14532), .op(n14564) );
  nand2_1 U11651 ( .ip1(n14496), .ip2(n14532), .op(n14500) );
  nand2_1 U11652 ( .ip1(n14482), .ip2(n14532), .op(n14489) );
  buf_2 U11653 ( .ip(n11999), .op(n13162) );
  nand2_4 U11654 ( .ip1(n14240), .ip2(n14030), .op(n14090) );
  buf_4 U11655 ( .ip(n14080), .op(n14404) );
  inv_2 U11656 ( .ip(n14090), .op(n14235) );
  nand2_2 U11657 ( .ip1(n14582), .ip2(n14581), .op(n19689) );
  nand2_1 U11658 ( .ip1(n14020), .ip2(n16525), .op(n14021) );
  nand2_1 U11659 ( .ip1(n14019), .ip2(n14018), .op(n14020) );
  buf_4 U11660 ( .ip(n14080), .op(n18024) );
  nand2_1 U11661 ( .ip1(n14489), .ip2(n14488), .op(n14490) );
  nand2_1 U11662 ( .ip1(n14477), .ip2(n14476), .op(n14491) );
  nand2_1 U11663 ( .ip1(n13575), .ip2(n13574), .op(n13579) );
  inv_2 U11664 ( .ip(n13166), .op(n16776) );
  inv_2 U11665 ( .ip(n19185), .op(n13166) );
  nand2_4 U11666 ( .ip1(n14308), .ip2(n10212), .op(n17433) );
  and2_2 U11667 ( .ip1(n14307), .ip2(n14306), .op(n10212) );
  nand2_2 U11668 ( .ip1(n11920), .ip2(n11919), .op(n21276) );
  or2_1 U11669 ( .ip1(n17399), .ip2(n11877), .op(n11920) );
  nand2_1 U11670 ( .ip1(imem_haddr[31]), .ip2(n21995), .op(n21987) );
  nand2_1 U11671 ( .ip1(n10205), .ip2(n20690), .op(n14286) );
  nand2_1 U11672 ( .ip1(n20690), .ip2(n20692), .op(n14297) );
  nand2_1 U11673 ( .ip1(n19894), .ip2(n14365), .op(n14370) );
  nand2_1 U11674 ( .ip1(n14120), .ip2(n14119), .op(n14078) );
  and2_2 U11675 ( .ip1(n21531), .ip2(n13753), .op(n10211) );
  nand2_1 U11676 ( .ip1(n12881), .ip2(n13315), .op(n17297) );
  nand2_1 U11677 ( .ip1(n11825), .ip2(n13315), .op(n11826) );
  nand2_2 U11678 ( .ip1(n13323), .ip2(n13322), .op(n13525) );
  nand2_1 U11679 ( .ip1(n10508), .ip2(n13315), .op(n10509) );
  or2_1 U11680 ( .ip1(n13315), .ip2(n11784), .op(n11827) );
  inv_2 U11681 ( .ip(n14090), .op(n14339) );
  nand2_2 U11682 ( .ip1(n12686), .ip2(n12685), .op(n17457) );
  nand2_4 U11683 ( .ip1(n10222), .ip2(n10454), .op(n13063) );
  xor2_2 U11684 ( .ip1(n17438), .ip2(n21994), .op(imem_haddr[2]) );
  nor2_1 U11685 ( .ip1(n14551), .ip2(n14547), .op(n10202) );
  and2_1 U11686 ( .ip1(n13785), .ip2(n10219), .op(n10203) );
  nand2_1 U11687 ( .ip1(n14392), .ip2(n14241), .op(n14030) );
  and2_1 U11688 ( .ip1(n13876), .ip2(n13875), .op(n10204) );
  and2_1 U11689 ( .ip1(n14579), .ip2(n14270), .op(n10205) );
  inv_2 U11690 ( .ip(n14339), .op(n14340) );
  inv_2 U11691 ( .ip(n14339), .op(n14413) );
  and2_1 U11692 ( .ip1(n14547), .ip2(n14552), .op(n10208) );
  and2_1 U11693 ( .ip1(n14195), .ip2(n14210), .op(n10213) );
  xor2_2 U11694 ( .ip1(n14390), .ip2(n14389), .op(imem_haddr[24]) );
  and2_1 U11695 ( .ip1(n14510), .ip2(n14507), .op(n10215) );
  and2_1 U11696 ( .ip1(n11952), .ip2(n11951), .op(n10216) );
  and2_1 U11697 ( .ip1(n14346), .ip2(n14345), .op(n10217) );
  nand2_1 U11698 ( .ip1(n13994), .ip2(n13858), .op(n18373) );
  inv_1 U11699 ( .ip(n11999), .op(n12184) );
  or2_1 U11700 ( .ip1(n10207), .ip2(n10184), .op(n10218) );
  and2_1 U11701 ( .ip1(n13784), .ip2(n13783), .op(n10219) );
  and2_1 U11702 ( .ip1(n11948), .ip2(n11947), .op(n10220) );
  and2_1 U11703 ( .ip1(n14565), .ip2(n14564), .op(n10221) );
  and2_1 U11704 ( .ip1(n10453), .ip2(n10452), .op(n10222) );
  and3_1 U11705 ( .ip1(n13610), .ip2(n13609), .ip3(n13608), .op(n10223) );
  nand2_1 U11706 ( .ip1(n14293), .ip2(n14294), .op(n20690) );
  and2_1 U11707 ( .ip1(n13900), .ip2(n13899), .op(n10224) );
  nor2_1 U11708 ( .ip1(n16533), .ip2(n13601), .op(n11945) );
  and2_1 U11709 ( .ip1(n13924), .ip2(n13921), .op(n10225) );
  and3_1 U11710 ( .ip1(n13931), .ip2(n13934), .ip3(n13935), .op(n10226) );
  and2_1 U11711 ( .ip1(n13883), .ip2(n13882), .op(n10227) );
  and2_1 U11712 ( .ip1(n13912), .ip2(n13911), .op(n10228) );
  nand2_1 U11713 ( .ip1(n12595), .ip2(n12594), .op(n12596) );
  and2_1 U11714 ( .ip1(n13704), .ip2(n13703), .op(n10229) );
  nand2_1 U11715 ( .ip1(n10181), .ip2(n17102), .op(n13899) );
  and2_1 U11716 ( .ip1(n13995), .ip2(n11936), .op(n10230) );
  inv_1 U11717 ( .ip(n13779), .op(n13983) );
  nand2_1 U11718 ( .ip1(n19069), .ip2(n10180), .op(n13779) );
  and2_1 U11719 ( .ip1(n12882), .ip2(n17296), .op(n10231) );
  and2_1 U11720 ( .ip1(n13980), .ip2(n13979), .op(n10232) );
  and2_1 U11721 ( .ip1(n16525), .ip2(n13748), .op(n10233) );
  and2_1 U11722 ( .ip1(n10190), .ip2(n16557), .op(n13643) );
  nor2_1 U11723 ( .ip1(n14445), .ip2(n14359), .op(n10234) );
  or2_1 U11724 ( .ip1(n14497), .ip2(n14453), .op(n10235) );
  inv_1 U11725 ( .ip(n13960), .op(n12139) );
  or2_1 U11726 ( .ip1(n13669), .ip2(n13668), .op(n10236) );
  nand2_1 U11727 ( .ip1(n16446), .ip2(n17584), .op(n13933) );
  inv_1 U11728 ( .ip(n13962), .op(n13963) );
  inv_1 U11729 ( .ip(n14276), .op(n14274) );
  nor2_1 U11730 ( .ip1(n10178), .ip2(n16935), .op(n13981) );
  nand2_1 U11731 ( .ip1(n13268), .ip2(n13267), .op(n13721) );
  nand2_1 U11732 ( .ip1(n18920), .ip2(n10191), .op(n13977) );
  inv_1 U11733 ( .ip(n13977), .op(n13778) );
  nand2_1 U11734 ( .ip1(n10193), .ip2(n13537), .op(n13932) );
  inv_1 U11735 ( .ip(n13932), .op(n13915) );
  inv_1 U11736 ( .ip(n14030), .op(n14031) );
  and2_1 U11737 ( .ip1(n20041), .ip2(n20037), .op(n10237) );
  nand3_1 U11738 ( .ip1(n14377), .ip2(n14381), .ip3(n14330), .op(n20037) );
  inv_1 U11739 ( .ip(n20037), .op(n20040) );
  nand2_1 U11740 ( .ip1(n14065), .ip2(n14064), .op(n14504) );
  inv_1 U11741 ( .ip(n14302), .op(n14589) );
  inv_1 U11742 ( .ip(n19687), .op(n14269) );
  inv_1 U11743 ( .ip(n14241), .op(n14029) );
  xor2_1 U11744 ( .ip1(n17517), .ip2(n20878), .op(n10239) );
  inv_1 U11745 ( .ip(n16445), .op(n16446) );
  inv_1 U11746 ( .ip(n18920), .op(n13600) );
  buf_1 U11747 ( .ip(n16913), .op(n20855) );
  inv_1 U11748 ( .ip(n16913), .op(n13613) );
  inv_1 U11749 ( .ip(n13754), .op(n13578) );
  nand2_1 U11840 ( .ip1(ext_interrupts[16]), .ip2(\pipeline/csr/mie [24]), 
        .op(n10241) );
  nand2_1 U11841 ( .ip1(\pipeline/csr/mie [25]), .ip2(ext_interrupts[17]), 
        .op(n10240) );
  nand2_1 U11842 ( .ip1(n10241), .ip2(n10240), .op(n10242) );
  not_ab_or_c_or_d U11843 ( .ip1(ext_interrupts[21]), .ip2(
        \pipeline/csr/mie [29]), .ip3(n10179), .ip4(n10242), .op(n10251) );
  nand2_1 U11844 ( .ip1(ext_interrupts[18]), .ip2(\pipeline/csr/mie [26]), 
        .op(n10244) );
  nand2_1 U11845 ( .ip1(ext_interrupts[4]), .ip2(\pipeline/csr/mie [12]), .op(
        n10243) );
  nand2_1 U11846 ( .ip1(n10244), .ip2(n10243), .op(n10246) );
  not_ab_or_c_or_d U11847 ( .ip1(\pipeline/csr/mie [30]), .ip2(
        ext_interrupts[22]), .ip3(n10246), .ip4(n10245), .op(n10250) );
  xor2_1 U11848 ( .ip1(\pipeline/prv [0]), .ip2(\pipeline/prv [1]), .op(n10248) );
  and2_1 U11849 ( .ip1(\pipeline/csr/mip_3 ), .ip2(\pipeline/csr/mie [3]), 
        .op(n10247) );
  not_ab_or_c_or_d U11850 ( .ip1(\pipeline/csr/mie [7]), .ip2(
        \pipeline/csr/mip[7] ), .ip3(n10248), .ip4(n10247), .op(n10249) );
  nand3_1 U11851 ( .ip1(n10251), .ip2(n10250), .ip3(n10249), .op(n10275) );
  nand2_1 U11852 ( .ip1(ext_interrupts[14]), .ip2(\pipeline/csr/mie [22]), 
        .op(n10255) );
  nand2_1 U11853 ( .ip1(ext_interrupts[12]), .ip2(\pipeline/csr/mie [20]), 
        .op(n10254) );
  nand2_1 U11854 ( .ip1(ext_interrupts[11]), .ip2(\pipeline/csr/mie [19]), 
        .op(n10253) );
  nand2_1 U11855 ( .ip1(ext_interrupts[15]), .ip2(\pipeline/csr/mie [23]), 
        .op(n10252) );
  nand4_1 U11856 ( .ip1(n10255), .ip2(n10254), .ip3(n10253), .ip4(n10252), 
        .op(n10261) );
  nand2_1 U11857 ( .ip1(ext_interrupts[9]), .ip2(\pipeline/csr/mie [17]), .op(
        n10259) );
  nand2_1 U11858 ( .ip1(ext_interrupts[7]), .ip2(\pipeline/csr/mie [15]), .op(
        n10258) );
  nand2_1 U11859 ( .ip1(ext_interrupts[10]), .ip2(\pipeline/csr/mie [18]), 
        .op(n10257) );
  nand2_1 U11860 ( .ip1(ext_interrupts[13]), .ip2(\pipeline/csr/mie [21]), 
        .op(n10256) );
  nand4_1 U11861 ( .ip1(n10259), .ip2(n10258), .ip3(n10257), .ip4(n10256), 
        .op(n10260) );
  nor2_1 U11862 ( .ip1(n10261), .ip2(n10260), .op(n10273) );
  nand2_1 U11863 ( .ip1(ext_interrupts[3]), .ip2(\pipeline/csr/mie [11]), .op(
        n10265) );
  nand2_1 U11864 ( .ip1(ext_interrupts[1]), .ip2(\pipeline/csr/mie [9]), .op(
        n10264) );
  nand2_1 U11865 ( .ip1(\pipeline/csr/mie [8]), .ip2(ext_interrupts[0]), .op(
        n10263) );
  nand2_1 U11866 ( .ip1(ext_interrupts[23]), .ip2(\pipeline/csr/mie [31]), 
        .op(n10262) );
  nand4_1 U11867 ( .ip1(n10265), .ip2(n10264), .ip3(n10263), .ip4(n10262), 
        .op(n10271) );
  nand2_1 U11868 ( .ip1(ext_interrupts[5]), .ip2(\pipeline/csr/mie [13]), .op(
        n10269) );
  nand2_1 U11869 ( .ip1(\pipeline/csr/mie [14]), .ip2(ext_interrupts[6]), .op(
        n10268) );
  nand2_1 U11870 ( .ip1(\pipeline/csr/mie [16]), .ip2(ext_interrupts[8]), .op(
        n10267) );
  nand2_1 U11871 ( .ip1(\pipeline/csr/mie [10]), .ip2(ext_interrupts[2]), .op(
        n10266) );
  nand4_1 U11872 ( .ip1(n10269), .ip2(n10268), .ip3(n10267), .ip4(n10266), 
        .op(n10270) );
  nor2_1 U11873 ( .ip1(n10271), .ip2(n10270), .op(n10272) );
  nand2_1 U11874 ( .ip1(n10273), .ip2(n10272), .op(n10274) );
  nor2_2 U11875 ( .ip1(n10275), .ip2(n10274), .op(n10289) );
  inv_1 U11876 ( .ip(n10289), .op(n10278) );
  inv_1 U11877 ( .ip(\pipeline/csr/priv_stack_0 ), .op(n10276) );
  nand3_1 U11878 ( .ip1(\pipeline/prv [1]), .ip2(\pipeline/prv [0]), .ip3(
        n10276), .op(n10277) );
  nand2_1 U11879 ( .ip1(n10278), .ip2(n10277), .op(n16055) );
  inv_1 U11880 ( .ip(n10294), .op(n21082) );
  inv_1 U11881 ( .ip(n10364), .op(n14034) );
  nor4_1 U11882 ( .ip1(ext_interrupts[22]), .ip2(ext_interrupts[20]), .ip3(
        ext_interrupts[18]), .ip4(ext_interrupts[4]), .op(n10282) );
  nor4_1 U11883 ( .ip1(ext_interrupts[21]), .ip2(ext_interrupts[19]), .ip3(
        ext_interrupts[16]), .ip4(ext_interrupts[17]), .op(n10281) );
  inv_1 U11884 ( .ip(\pipeline/ctrl/wfi_unkilled_WB ), .op(n10279) );
  nor4_1 U11885 ( .ip1(\pipeline/csr/mip[7] ), .ip2(\pipeline/csr/mip_3 ), 
        .ip3(\pipeline/ctrl/prev_killed_WB ), .ip4(n10279), .op(n10280) );
  nand3_1 U11886 ( .ip1(n10282), .ip2(n10281), .ip3(n10280), .op(n10288) );
  nor4_2 U11887 ( .ip1(ext_interrupts[14]), .ip2(ext_interrupts[15]), .ip3(
        ext_interrupts[13]), .ip4(ext_interrupts[11]), .op(n10286) );
  nor4_2 U11888 ( .ip1(ext_interrupts[12]), .ip2(ext_interrupts[9]), .ip3(
        ext_interrupts[10]), .ip4(ext_interrupts[7]), .op(n10285) );
  nor4_2 U11889 ( .ip1(ext_interrupts[8]), .ip2(ext_interrupts[6]), .ip3(
        ext_interrupts[5]), .ip4(ext_interrupts[2]), .op(n10284) );
  nor4_2 U11890 ( .ip1(ext_interrupts[3]), .ip2(ext_interrupts[0]), .ip3(
        ext_interrupts[23]), .ip4(ext_interrupts[1]), .op(n10283) );
  nand4_1 U11891 ( .ip1(n10286), .ip2(n10285), .ip3(n10284), .ip4(n10283), 
        .op(n10287) );
  nor2_2 U11892 ( .ip1(n10288), .ip2(n10287), .op(n10366) );
  inv_1 U11893 ( .ip(dmem_hready), .op(n10290) );
  nand2_1 U11894 ( .ip1(n10290), .ip2(\pipeline/ctrl/dmem_en_WB ), .op(n10293)
         );
  nand2_1 U11895 ( .ip1(\pipeline/md/state [0]), .ip2(\pipeline/md/state [1]), 
        .op(n10291) );
  nand2_1 U11896 ( .ip1(\pipeline/ctrl/uses_md_WB ), .ip2(n10291), .op(n10292)
         );
  nand2_1 U11897 ( .ip1(n10293), .ip2(n10292), .op(n10450) );
  nand2_1 U11898 ( .ip1(n10294), .ip2(\pipeline/ctrl/wr_reg_unkilled_WB ), 
        .op(n10449) );
  nor2_1 U11899 ( .ip1(n10450), .ip2(n10449), .op(n10443) );
  nand2_1 U11900 ( .ip1(n10454), .ip2(n10443), .op(n10295) );
  inv_1 U11901 ( .ip(n10295), .op(n17907) );
  inv_1 U11902 ( .ip(\pipeline/inst_DX [18]), .op(n15821) );
  xor2_1 U11903 ( .ip1(\pipeline/reg_to_wr_WB [3]), .ip2(n15821), .op(n10438)
         );
  inv_1 U11904 ( .ip(n10438), .op(n10298) );
  xor2_1 U11905 ( .ip1(\pipeline/inst_DX [15]), .ip2(
        \pipeline/reg_to_wr_WB [0]), .op(n10436) );
  xor2_1 U11906 ( .ip1(\pipeline/inst_DX [17]), .ip2(
        \pipeline/reg_to_wr_WB [2]), .op(n10435) );
  or2_1 U11907 ( .ip1(\pipeline/inst_DX [17]), .ip2(\pipeline/inst_DX [19]), 
        .op(n10377) );
  nor2_1 U11908 ( .ip1(\pipeline/inst_DX [18]), .ip2(n10377), .op(n10381) );
  nor2_1 U11909 ( .ip1(\pipeline/inst_DX [16]), .ip2(\pipeline/inst_DX [15]), 
        .op(n10376) );
  nand2_1 U11910 ( .ip1(n10381), .ip2(n10376), .op(n15311) );
  inv_1 U11911 ( .ip(\pipeline/reg_to_wr_WB [4]), .op(n17906) );
  xor2_1 U11912 ( .ip1(\pipeline/inst_DX [19]), .ip2(n17906), .op(n10437) );
  xor2_1 U11913 ( .ip1(\pipeline/inst_DX [16]), .ip2(
        \pipeline/reg_to_wr_WB [1]), .op(n10434) );
  inv_1 U11914 ( .ip(n10434), .op(n10296) );
  nand3_1 U11915 ( .ip1(n15311), .ip2(n10437), .ip3(n10296), .op(n10297) );
  nand2_1 U11916 ( .ip1(\pipeline/inst_DX [4]), .ip2(\pipeline/inst_DX [2]), 
        .op(n10299) );
  nand2_1 U11917 ( .ip1(\pipeline/inst_DX [5]), .ip2(n10299), .op(n10303) );
  inv_1 U11918 ( .ip(\pipeline/inst_DX [3]), .op(n10372) );
  nor2_1 U11919 ( .ip1(\pipeline/inst_DX [5]), .ip2(n10372), .op(n10306) );
  inv_1 U11920 ( .ip(\pipeline/inst_DX [4]), .op(n10307) );
  nand2_1 U11921 ( .ip1(\pipeline/inst_DX [2]), .ip2(n10307), .op(n10304) );
  nor3_1 U11922 ( .ip1(\pipeline/inst_DX [6]), .ip2(n10306), .ip3(n10304), 
        .op(n10302) );
  nand2_1 U11923 ( .ip1(\pipeline/inst_DX [0]), .ip2(\pipeline/inst_DX [1]), 
        .op(n16483) );
  inv_1 U11924 ( .ip(n16483), .op(n17786) );
  nand2_1 U11925 ( .ip1(\pipeline/inst_DX [3]), .ip2(n10304), .op(n10300) );
  nand2_1 U11926 ( .ip1(n17786), .ip2(n10300), .op(n10301) );
  not_ab_or_c_or_d U11927 ( .ip1(\pipeline/inst_DX [6]), .ip2(n10303), .ip3(
        n10302), .ip4(n10301), .op(n10347) );
  inv_1 U11928 ( .ip(\pipeline/inst_DX [5]), .op(n17784) );
  nor2_1 U11929 ( .ip1(\pipeline/inst_DX [2]), .ip2(n17784), .op(n10313) );
  inv_1 U11930 ( .ip(n10313), .op(n10332) );
  inv_1 U11931 ( .ip(\pipeline/inst_DX [6]), .op(n10305) );
  nor3_1 U11932 ( .ip1(\pipeline/inst_DX [3]), .ip2(n10332), .ip3(n10305), 
        .op(n10308) );
  nand2_1 U11933 ( .ip1(n10308), .ip2(\pipeline/inst_DX [4]), .op(n15310) );
  inv_1 U11934 ( .ip(n10304), .op(n10311) );
  nand3_1 U11935 ( .ip1(n10311), .ip2(n10306), .ip3(n10305), .op(n10330) );
  or2_1 U11936 ( .ip1(\pipeline/inst_DX [3]), .ip2(\pipeline/inst_DX [6]), 
        .op(n10309) );
  nor3_1 U11937 ( .ip1(\pipeline/inst_DX [2]), .ip2(\pipeline/inst_DX [4]), 
        .ip3(n10309), .op(n17785) );
  inv_1 U11938 ( .ip(n17785), .op(n17740) );
  nand2_1 U11939 ( .ip1(n10308), .ip2(n10307), .op(n16479) );
  inv_1 U11940 ( .ip(n10309), .op(n10310) );
  nand2_1 U11941 ( .ip1(\pipeline/inst_DX [4]), .ip2(n10310), .op(n17886) );
  or2_1 U11942 ( .ip1(\pipeline/inst_DX [2]), .ip2(n17886), .op(n16477) );
  nand2_1 U11943 ( .ip1(n16479), .ip2(n16477), .op(n13576) );
  nor2_1 U11944 ( .ip1(n10314), .ip2(n13576), .op(n10511) );
  nand2_1 U11945 ( .ip1(\pipeline/inst_DX [6]), .ip2(n10311), .op(n10316) );
  inv_1 U11946 ( .ip(n10316), .op(n13210) );
  nand2_1 U11947 ( .ip1(n13210), .ip2(n10372), .op(n10344) );
  nand2_1 U11948 ( .ip1(n10511), .ip2(n10344), .op(n10441) );
  nand3_1 U11949 ( .ip1(n17907), .ip2(n10312), .ip3(n10441), .op(n10325) );
  nand3_1 U11950 ( .ip1(\pipeline/inst_DX [5]), .ip2(n17786), .ip3(n17785), 
        .op(n13443) );
  nor2_1 U11951 ( .ip1(n10313), .ip2(n17886), .op(n10315) );
  nor2_1 U11952 ( .ip1(n10315), .ip2(n10314), .op(n13209) );
  nand2_1 U11953 ( .ip1(n13209), .ip2(n10316), .op(n12091) );
  nor2_1 U11954 ( .ip1(\pipeline/inst_DX [24]), .ip2(\pipeline/inst_DX [22]), 
        .op(n10464) );
  inv_1 U11955 ( .ip(\pipeline/inst_DX [23]), .op(n13117) );
  nand2_1 U11956 ( .ip1(n10464), .ip2(n13117), .op(n15340) );
  or2_1 U11957 ( .ip1(\pipeline/inst_DX [21]), .ip2(\pipeline/inst_DX [20]), 
        .op(n22094) );
  nor2_1 U11958 ( .ip1(n15340), .ip2(n22094), .op(n22119) );
  xor2_1 U11959 ( .ip1(\pipeline/inst_DX [23]), .ip2(
        \pipeline/reg_to_wr_WB [3]), .op(n10319) );
  xor2_1 U11960 ( .ip1(\pipeline/inst_DX [21]), .ip2(
        \pipeline/reg_to_wr_WB [1]), .op(n10318) );
  xor2_1 U11961 ( .ip1(\pipeline/inst_DX [22]), .ip2(
        \pipeline/reg_to_wr_WB [2]), .op(n10317) );
  nor3_1 U11962 ( .ip1(n10319), .ip2(n10318), .ip3(n10317), .op(n10322) );
  xor2_1 U11963 ( .ip1(\pipeline/inst_DX [24]), .ip2(n17906), .op(n10321) );
  inv_1 U11964 ( .ip(\pipeline/reg_to_wr_WB [0]), .op(n17908) );
  xor2_1 U11965 ( .ip1(\pipeline/inst_DX [20]), .ip2(n17908), .op(n10320) );
  nand3_1 U11966 ( .ip1(n10322), .ip2(n10321), .ip3(n10320), .op(n10323) );
  not_ab_or_c_or_d U11967 ( .ip1(n13443), .ip2(n12091), .ip3(n22119), .ip4(
        n10323), .op(n10452) );
  nand2_1 U11968 ( .ip1(n17907), .ip2(n10452), .op(n10324) );
  nand2_1 U11969 ( .ip1(n10325), .ip2(n10324), .op(n10327) );
  inv_1 U11970 ( .ip(\pipeline/ctrl/dmem_en_WB ), .op(n10326) );
  nor2_1 U11971 ( .ip1(\pipeline/ctrl/store_in_WB ), .ip2(n10326), .op(n10451)
         );
  nand2_1 U11972 ( .ip1(n10327), .ip2(n10451), .op(n10336) );
  or3_1 U11973 ( .ip1(\pipeline/inst_DX [9]), .ip2(\pipeline/inst_DX [7]), 
        .ip3(\pipeline/inst_DX [8]), .op(n10328) );
  nor4_1 U11974 ( .ip1(\pipeline/inst_DX [11]), .ip2(\pipeline/inst_DX [10]), 
        .ip3(n15311), .ip4(n10328), .op(n10353) );
  nor2_1 U11975 ( .ip1(\pipeline/inst_DX [26]), .ip2(\pipeline/inst_DX [25]), 
        .op(n15330) );
  nor3_1 U11976 ( .ip1(\pipeline/imm[31] ), .ip2(\pipeline/inst_DX [30]), 
        .ip3(\pipeline/inst_DX [29]), .op(n10354) );
  inv_1 U11977 ( .ip(n15340), .op(n22112) );
  inv_1 U11978 ( .ip(\pipeline/inst_DX [27]), .op(n15339) );
  nor2_1 U11979 ( .ip1(\pipeline/dmem_type[2] ), .ip2(dmem_hsize[1]), .op(
        n16478) );
  inv_1 U11980 ( .ip(n16478), .op(n10341) );
  nor4_1 U11981 ( .ip1(\pipeline/inst_DX [28]), .ip2(n10343), .ip3(n10341), 
        .ip4(n22094), .op(n10329) );
  nand2_1 U11982 ( .ip1(n10353), .ip2(n10329), .op(n10356) );
  inv_1 U11983 ( .ip(n10330), .op(n10357) );
  nand4_1 U11984 ( .ip1(n10357), .ip2(n17786), .ip3(dmem_hsize[0]), .ip4(
        \pipeline/ctrl/store_in_WB ), .op(n10331) );
  nor2_1 U11985 ( .ip1(n10356), .ip2(n10331), .op(n17744) );
  nor2_1 U11986 ( .ip1(\pipeline/md/state [0]), .ip2(\pipeline/md/state [1]), 
        .op(n14771) );
  nor2_1 U11987 ( .ip1(n10332), .ip2(n17886), .op(n13582) );
  inv_1 U11988 ( .ip(\pipeline/inst_DX [26]), .op(n11367) );
  nand2_1 U11989 ( .ip1(\pipeline/inst_DX [25]), .ip2(n11367), .op(n15332) );
  nor4_1 U11990 ( .ip1(\pipeline/inst_DX [27]), .ip2(\pipeline/inst_DX [28]), 
        .ip3(n16483), .ip4(n15332), .op(n10333) );
  nand3_1 U11991 ( .ip1(n10354), .ip2(n13582), .ip3(n10333), .op(n17788) );
  nor2_1 U11992 ( .ip1(n14771), .ip2(n17788), .op(n10334) );
  nor2_1 U11993 ( .ip1(n17744), .ip2(n10334), .op(n10335) );
  nand2_1 U11994 ( .ip1(n10336), .ip2(n10335), .op(n10365) );
  inv_1 U11995 ( .ip(dmem_hsize[0]), .op(n15312) );
  inv_1 U11996 ( .ip(dmem_hsize[1]), .op(n15352) );
  nand2_1 U11997 ( .ip1(n15312), .ip2(n15352), .op(n22090) );
  nor2_1 U11998 ( .ip1(n15310), .ip2(n22090), .op(n10361) );
  inv_1 U11999 ( .ip(\pipeline/inst_DX [28]), .op(n22120) );
  nor2_1 U12000 ( .ip1(\pipeline/prv [0]), .ip2(\pipeline/prv [1]), .op(n10337) );
  nor2_1 U12001 ( .ip1(n10337), .ip2(n22094), .op(n14025) );
  inv_1 U12002 ( .ip(\pipeline/inst_DX [20]), .op(n11079) );
  nand2_1 U12003 ( .ip1(\pipeline/inst_DX [21]), .ip2(n11079), .op(n17317) );
  inv_1 U12004 ( .ip(n17317), .op(n17778) );
  nor3_1 U12005 ( .ip1(n14025), .ip2(n17778), .ip3(n22120), .op(n10338) );
  not_ab_or_c_or_d U12006 ( .ip1(\pipeline/inst_DX [21]), .ip2(n22120), .ip3(
        n10338), .ip4(n10343), .op(n10339) );
  inv_1 U12007 ( .ip(n10353), .op(n10342) );
  nor2_1 U12008 ( .ip1(n10339), .ip2(n10342), .op(n10340) );
  or2_1 U12009 ( .ip1(\pipeline/dmem_type[2] ), .ip2(n10340), .op(n10360) );
  nor2_1 U12010 ( .ip1(dmem_hsize[0]), .ip2(n10341), .op(n14596) );
  inv_1 U12011 ( .ip(n14596), .op(n17883) );
  nand2_1 U12012 ( .ip1(n17779), .ip2(n22120), .op(n10362) );
  inv_1 U12013 ( .ip(\pipeline/inst_DX [21]), .op(n13319) );
  nand2_1 U12014 ( .ip1(\pipeline/inst_DX [20]), .ip2(n13319), .op(n15315) );
  nor2_1 U12015 ( .ip1(n10362), .ip2(n15315), .op(n18388) );
  inv_1 U12016 ( .ip(\pipeline/dmem_type[2] ), .op(n17765) );
  nand2_1 U12017 ( .ip1(dmem_hsize[1]), .ip2(n17765), .op(n13577) );
  inv_1 U12018 ( .ip(n13577), .op(n16480) );
  inv_1 U12019 ( .ip(n16479), .op(n10352) );
  inv_1 U12020 ( .ip(n10344), .op(n10345) );
  nand2_1 U12021 ( .ip1(n10345), .ip2(n17883), .op(n10346) );
  nand2_1 U12022 ( .ip1(n10347), .ip2(n10346), .op(n10351) );
  nand3_1 U12023 ( .ip1(\pipeline/imm[31] ), .ip2(\pipeline/inst_DX [30]), 
        .ip3(\pipeline/csr/system_wen ), .op(n10349) );
  nor2_1 U12024 ( .ip1(\pipeline/csr/N2385 ), .ip2(\pipeline/csr/N2387 ), .op(
        n10348) );
  nand2_1 U12025 ( .ip1(n10349), .ip2(n10348), .op(n10350) );
  not_ab_or_c_or_d U12026 ( .ip1(n16480), .ip2(n10352), .ip3(n10351), .ip4(
        n10350), .op(n10359) );
  nand3_1 U12027 ( .ip1(n10357), .ip2(n10356), .ip3(n10355), .op(n10358) );
  nand2_1 U12028 ( .ip1(n10359), .ip2(n10358), .op(n18386) );
  not_ab_or_c_or_d U12029 ( .ip1(n10361), .ip2(n10360), .ip3(n18388), .ip4(
        n18386), .op(n21097) );
  inv_1 U12030 ( .ip(n10362), .op(n21095) );
  nor2_1 U12031 ( .ip1(n21095), .ip2(\pipeline/ctrl/had_ex_DX ), .op(n10363)
         );
  nand2_1 U12032 ( .ip1(n21097), .ip2(n10363), .op(n22046) );
  nand2_1 U12033 ( .ip1(n10365), .ip2(n17674), .op(n10369) );
  nand2_1 U12034 ( .ip1(n16055), .ip2(n10366), .op(n10368) );
  inv_1 U12035 ( .ip(n10450), .op(n10367) );
  nand2_1 U12036 ( .ip1(n10368), .ip2(n10367), .op(n17320) );
  nand2_1 U12037 ( .ip1(n17320), .ip2(n20972), .op(n17741) );
  and2_1 U12038 ( .ip1(n10369), .ip2(n17741), .op(n17816) );
  inv_1 U12039 ( .ip(n17816), .op(n17804) );
  nand2_1 U12040 ( .ip1(n17804), .ip2(imem_hready), .op(n10370) );
  inv_1 U12041 ( .ip(\pipeline/ctrl/replay_IF ), .op(n17673) );
  and2_1 U12042 ( .ip1(n10370), .ip2(n17673), .op(n14032) );
  inv_1 U12043 ( .ip(n14032), .op(n10371) );
  nor2_1 U12044 ( .ip1(n10364), .ip2(n10371), .op(n14169) );
  inv_1 U12045 ( .ip(n17819), .op(n17891) );
  and2_1 U12046 ( .ip1(n17891), .ip2(n13210), .op(n17888) );
  inv_1 U12047 ( .ip(\pipeline/wb_src_sel_WB [1]), .op(n17895) );
  nor2_1 U12048 ( .ip1(\pipeline/wb_src_sel_WB [0]), .ip2(n17895), .op(n13368)
         );
  nand2_1 U12049 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [19]), .op(n10375) );
  nand2_1 U12050 ( .ip1(\pipeline/alu_out_WB [19]), .ip2(n17895), .op(n10374)
         );
  nand2_1 U12051 ( .ip1(\pipeline/wb_src_sel_WB [1]), .ip2(
        \pipeline/wb_src_sel_WB [0]), .op(n13217) );
  inv_1 U12052 ( .ip(n13217), .op(n13369) );
  nand2_1 U12053 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [19]), .op(
        n10373) );
  nand3_1 U12054 ( .ip1(n10375), .ip2(n10374), .ip3(n10373), .op(n18579) );
  inv_1 U12055 ( .ip(n10376), .op(n10421) );
  inv_1 U12056 ( .ip(\pipeline/inst_DX [17]), .op(n15782) );
  nor2_1 U12057 ( .ip1(n15782), .ip2(n15821), .op(n10411) );
  nand2_1 U12058 ( .ip1(\pipeline/inst_DX [19]), .ip2(n10411), .op(n10419) );
  nor2_1 U12059 ( .ip1(n10421), .ip2(n10419), .op(n13462) );
  inv_1 U12060 ( .ip(n10377), .op(n10378) );
  nand2_1 U12061 ( .ip1(n10378), .ip2(\pipeline/inst_DX [18]), .op(n10404) );
  nor2_1 U12062 ( .ip1(n10421), .ip2(n10404), .op(n13448) );
  nand2_1 U12063 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][19] ), .op(
        n10380) );
  inv_1 U12064 ( .ip(\pipeline/inst_DX [15]), .op(n16028) );
  nand2_1 U12065 ( .ip1(\pipeline/inst_DX [16]), .ip2(n16028), .op(n10418) );
  nor2_1 U12066 ( .ip1(n10404), .ip2(n10418), .op(n13449) );
  nand2_1 U12067 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][19] ), .op(
        n10379) );
  nand2_1 U12068 ( .ip1(n10380), .ip2(n10379), .op(n10387) );
  inv_1 U12069 ( .ip(\pipeline/inst_DX [16]), .op(n15833) );
  nand2_1 U12070 ( .ip1(\pipeline/inst_DX [15]), .ip2(n15833), .op(n10417) );
  nand3_1 U12071 ( .ip1(\pipeline/inst_DX [19]), .ip2(\pipeline/inst_DX [17]), 
        .ip3(n15821), .op(n10410) );
  nor2_1 U12072 ( .ip1(n10417), .ip2(n10410), .op(n13452) );
  nand2_1 U12073 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][19] ), .op(
        n10385) );
  inv_1 U12074 ( .ip(\pipeline/inst_DX [19]), .op(n15660) );
  nor2_1 U12075 ( .ip1(\pipeline/inst_DX [17]), .ip2(n15660), .op(n10388) );
  nand2_1 U12076 ( .ip1(n10388), .ip2(n15821), .op(n10405) );
  nor2_1 U12077 ( .ip1(n10417), .ip2(n10405), .op(n13453) );
  nand2_1 U12078 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][19] ), .op(
        n10384) );
  nand2_1 U12079 ( .ip1(\pipeline/inst_DX [16]), .ip2(\pipeline/inst_DX [15]), 
        .op(n10412) );
  nand3_1 U12080 ( .ip1(\pipeline/inst_DX [17]), .ip2(n15821), .ip3(n15660), 
        .op(n10399) );
  nor2_1 U12081 ( .ip1(n10412), .ip2(n10399), .op(n13454) );
  nand2_1 U12082 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][19] ), .op(
        n10383) );
  inv_1 U12083 ( .ip(n10381), .op(n10398) );
  nor2_1 U12084 ( .ip1(n10398), .ip2(n10417), .op(n13455) );
  nand2_1 U12085 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][19] ), .op(
        n10382) );
  not_ab_or_c_or_d U12086 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][19] ), .ip3(n10387), .ip4(n10386), .op(n10433) );
  nand2_1 U12087 ( .ip1(\pipeline/inst_DX [18]), .ip2(n10388), .op(n10397) );
  nor2_1 U12088 ( .ip1(n10412), .ip2(n10397), .op(n13463) );
  nand2_1 U12089 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][19] ), .op(
        n10392) );
  nor2_1 U12090 ( .ip1(n10404), .ip2(n10417), .op(n13464) );
  nand2_1 U12091 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][19] ), .op(
        n10391) );
  nor2_1 U12092 ( .ip1(n10398), .ip2(n10418), .op(n13465) );
  nand2_1 U12093 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][19] ), .op(
        n10390) );
  nor2_1 U12094 ( .ip1(n10418), .ip2(n10397), .op(n13466) );
  nand2_1 U12095 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][19] ), .op(
        n10389) );
  and4_1 U12096 ( .ip1(n10392), .ip2(n10391), .ip3(n10390), .ip4(n10389), .op(
        n10432) );
  nor2_1 U12097 ( .ip1(n10421), .ip2(n10405), .op(n13471) );
  nand2_1 U12098 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][19] ), .op(
        n10396) );
  nor2_1 U12099 ( .ip1(n10421), .ip2(n10399), .op(n13472) );
  nand2_1 U12100 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][19] ), .op(
        n10395) );
  nor2_1 U12101 ( .ip1(n10421), .ip2(n10397), .op(n13473) );
  nand2_1 U12102 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][19] ), .op(
        n10394) );
  nor2_1 U12103 ( .ip1(n10421), .ip2(n10410), .op(n13474) );
  nand2_1 U12104 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][19] ), .op(
        n10393) );
  and4_1 U12105 ( .ip1(n10396), .ip2(n10395), .ip3(n10394), .ip4(n10393), .op(
        n10431) );
  nor2_1 U12106 ( .ip1(n10417), .ip2(n10397), .op(n13479) );
  nand2_1 U12107 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][19] ), .op(
        n10403) );
  nor2_1 U12108 ( .ip1(n10398), .ip2(n10412), .op(n13480) );
  nand2_1 U12109 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][19] ), .op(
        n10402) );
  nor2_1 U12110 ( .ip1(n10418), .ip2(n10399), .op(n13481) );
  nand2_1 U12111 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][19] ), .op(
        n10401) );
  nor2_1 U12112 ( .ip1(n10417), .ip2(n10399), .op(n13482) );
  nand2_1 U12113 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][19] ), .op(
        n10400) );
  nor2_1 U12114 ( .ip1(n10418), .ip2(n10405), .op(n13487) );
  nand2_1 U12115 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][19] ), .op(
        n10409) );
  nor2_1 U12116 ( .ip1(n10410), .ip2(n10412), .op(n13488) );
  nand2_1 U12117 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][19] ), .op(
        n10408) );
  nor2_1 U12118 ( .ip1(n10404), .ip2(n10412), .op(n13489) );
  nand2_1 U12119 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][19] ), .op(
        n10407) );
  nor2_1 U12120 ( .ip1(n10405), .ip2(n10412), .op(n13490) );
  nand2_1 U12121 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][19] ), .op(
        n10406) );
  nor2_1 U12122 ( .ip1(n10419), .ip2(n10417), .op(n13495) );
  nand2_1 U12123 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][19] ), .op(
        n10416) );
  nor2_1 U12124 ( .ip1(n10418), .ip2(n10410), .op(n13496) );
  nand2_1 U12125 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][19] ), .op(
        n10415) );
  nand2_1 U12126 ( .ip1(n10411), .ip2(n15660), .op(n10420) );
  nor2_1 U12127 ( .ip1(n10412), .ip2(n10420), .op(n13497) );
  nand2_1 U12128 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][19] ), .op(
        n10414) );
  nor2_1 U12129 ( .ip1(n10419), .ip2(n10412), .op(n13498) );
  nand2_1 U12130 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][19] ), .op(
        n10413) );
  nor2_1 U12131 ( .ip1(n10418), .ip2(n10420), .op(n13503) );
  nand2_1 U12132 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][19] ), .op(
        n10425) );
  nor2_1 U12133 ( .ip1(n10417), .ip2(n10420), .op(n13504) );
  nand2_1 U12134 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][19] ), .op(
        n10424) );
  nor2_1 U12135 ( .ip1(n10419), .ip2(n10418), .op(n13505) );
  nand2_1 U12136 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][19] ), .op(
        n10423) );
  nor2_1 U12137 ( .ip1(n10421), .ip2(n10420), .op(n13506) );
  nand2_1 U12138 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][19] ), .op(
        n10422) );
  and4_1 U12139 ( .ip1(n10439), .ip2(n15311), .ip3(n10438), .ip4(n10437), .op(
        n10440) );
  nand2_2 U12140 ( .ip1(n10454), .ip2(n10444), .op(n11999) );
  buf_2 U12141 ( .ip(n11999), .op(n13364) );
  mux2_1 U12142 ( .ip1(n18579), .ip2(n10445), .s(n10199), .op(n15628) );
  inv_1 U12143 ( .ip(n10511), .op(n13520) );
  nand2_1 U12144 ( .ip1(n15628), .ip2(n13520), .op(n10448) );
  nor2_1 U12145 ( .ip1(n13210), .ip2(n17784), .op(n10446) );
  nor2_1 U12146 ( .ip1(n10446), .ip2(n13520), .op(n13521) );
  nand2_1 U12147 ( .ip1(n13521), .ip2(\pipeline/PC_DX [19]), .op(n10447) );
  nand2_1 U12148 ( .ip1(n10448), .ip2(n10447), .op(n13666) );
  inv_1 U12149 ( .ip(n13666), .op(n13617) );
  inv_1 U12150 ( .ip(n10188), .op(n10517) );
  nor3_1 U12151 ( .ip1(n10451), .ip2(n10450), .ip3(n10449), .op(n10453) );
  buf_4 U12152 ( .ip(n13063), .op(n13441) );
  nand2_1 U12153 ( .ip1(\pipeline/inst_DX [22]), .ip2(\pipeline/inst_DX [23]), 
        .op(n10492) );
  or2_1 U12154 ( .ip1(\pipeline/inst_DX [24]), .ip2(n10492), .op(n10487) );
  nor2_1 U12155 ( .ip1(n17317), .ip2(n10487), .op(n13384) );
  inv_1 U12156 ( .ip(\pipeline/inst_DX [24]), .op(n12837) );
  nand3_1 U12157 ( .ip1(\pipeline/inst_DX [22]), .ip2(n13117), .ip3(n12837), 
        .op(n10486) );
  nor2_1 U12158 ( .ip1(n22094), .ip2(n10486), .op(n22097) );
  nand2_1 U12159 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][19] ), .op(
        n10457) );
  nor2_1 U12160 ( .ip1(n15340), .ip2(n15315), .op(n22109) );
  nand2_1 U12161 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][19] ), .op(
        n10456) );
  nand2_1 U12162 ( .ip1(n10457), .ip2(n10456), .op(n10463) );
  nor2_1 U12163 ( .ip1(n15340), .ip2(n17317), .op(n15338) );
  nand2_1 U12164 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][19] ), .op(
        n10461) );
  nor2_1 U12165 ( .ip1(\pipeline/inst_DX [22]), .ip2(n12837), .op(n10465) );
  nand2_1 U12166 ( .ip1(n10465), .ip2(n13117), .op(n10475) );
  nor2_1 U12167 ( .ip1(n22094), .ip2(n10475), .op(n13375) );
  nand2_1 U12168 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][19] ), .op(
        n10460) );
  nand2_1 U12169 ( .ip1(\pipeline/inst_DX [20]), .ip2(\pipeline/inst_DX [21]), 
        .op(n10494) );
  or2_1 U12170 ( .ip1(n15340), .ip2(n10494), .op(n15309) );
  inv_1 U12171 ( .ip(n15309), .op(n13376) );
  nand2_1 U12172 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][19] ), .op(
        n10459) );
  nand3_1 U12173 ( .ip1(\pipeline/inst_DX [22]), .ip2(\pipeline/inst_DX [24]), 
        .ip3(n13117), .op(n10481) );
  nor2_1 U12174 ( .ip1(n22094), .ip2(n10481), .op(n13377) );
  nand2_1 U12175 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][19] ), .op(
        n10458) );
  not_ab_or_c_or_d U12176 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][19] ), .ip3(n10463), .ip4(n10462), .op(n10507) );
  nand2_1 U12177 ( .ip1(n10464), .ip2(\pipeline/inst_DX [23]), .op(n10474) );
  nor2_1 U12178 ( .ip1(n15315), .ip2(n10474), .op(n13385) );
  nand2_1 U12179 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][19] ), .op(
        n10469) );
  nor2_1 U12180 ( .ip1(n15315), .ip2(n10481), .op(n13386) );
  nand2_1 U12181 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][19] ), .op(
        n10468) );
  nand2_1 U12182 ( .ip1(\pipeline/inst_DX [23]), .ip2(n10465), .op(n10480) );
  nor2_1 U12183 ( .ip1(n22094), .ip2(n10480), .op(n13387) );
  nand2_1 U12184 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][19] ), .op(
        n10467) );
  nor2_1 U12185 ( .ip1(n17317), .ip2(n10474), .op(n13388) );
  nand2_1 U12186 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][19] ), .op(
        n10466) );
  and4_1 U12187 ( .ip1(n10469), .ip2(n10468), .ip3(n10467), .ip4(n10466), .op(
        n10506) );
  nor2_1 U12188 ( .ip1(n10486), .ip2(n10494), .op(n13393) );
  nand2_1 U12189 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][19] ), .op(
        n10473) );
  nor2_1 U12190 ( .ip1(n22094), .ip2(n10474), .op(n13394) );
  nand2_1 U12191 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][19] ), .op(
        n10472) );
  nor2_1 U12192 ( .ip1(n10494), .ip2(n10481), .op(n13395) );
  nand2_1 U12193 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][19] ), .op(
        n10471) );
  nor2_1 U12194 ( .ip1(n15315), .ip2(n10475), .op(n13396) );
  nand2_1 U12195 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][19] ), .op(
        n10470) );
  and4_1 U12196 ( .ip1(n10473), .ip2(n10472), .ip3(n10471), .ip4(n10470), .op(
        n10505) );
  nor2_1 U12197 ( .ip1(n10494), .ip2(n10474), .op(n13401) );
  nand2_1 U12198 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][19] ), .op(
        n10479) );
  nor2_1 U12199 ( .ip1(n15315), .ip2(n10480), .op(n13402) );
  nand2_1 U12200 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][19] ), .op(
        n10478) );
  nor2_1 U12201 ( .ip1(n17317), .ip2(n10475), .op(n13403) );
  nand2_1 U12202 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][19] ), .op(
        n10477) );
  nor2_1 U12203 ( .ip1(n10475), .ip2(n10494), .op(n13404) );
  nand2_1 U12204 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][19] ), .op(
        n10476) );
  nor2_1 U12205 ( .ip1(n17317), .ip2(n10486), .op(n13409) );
  nand2_1 U12206 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][19] ), .op(
        n10485) );
  nor2_1 U12207 ( .ip1(n10494), .ip2(n10480), .op(n13410) );
  nand2_1 U12208 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][19] ), .op(
        n10484) );
  nor2_1 U12209 ( .ip1(n17317), .ip2(n10480), .op(n13411) );
  nand2_1 U12210 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][19] ), .op(
        n10483) );
  nor2_1 U12211 ( .ip1(n17317), .ip2(n10481), .op(n13412) );
  nand2_1 U12212 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][19] ), .op(
        n10482) );
  nor2_1 U12213 ( .ip1(n10487), .ip2(n10494), .op(n13417) );
  nand2_1 U12214 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][19] ), .op(
        n10491) );
  nor2_1 U12215 ( .ip1(n15315), .ip2(n10486), .op(n13418) );
  nand2_1 U12216 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][19] ), .op(
        n10490) );
  nor2_1 U12217 ( .ip1(n22094), .ip2(n10487), .op(n13419) );
  nand2_1 U12218 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][19] ), .op(
        n10489) );
  nor2_1 U12219 ( .ip1(n15315), .ip2(n10487), .op(n13420) );
  nand2_1 U12220 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][19] ), .op(
        n10488) );
  inv_1 U12221 ( .ip(n10492), .op(n10493) );
  nand2_1 U12222 ( .ip1(n10493), .ip2(\pipeline/inst_DX [24]), .op(n10495) );
  nor2_1 U12223 ( .ip1(n17317), .ip2(n10495), .op(n13425) );
  nand2_1 U12224 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][19] ), .op(
        n10499) );
  nor2_1 U12225 ( .ip1(n22094), .ip2(n10495), .op(n13426) );
  nand2_1 U12226 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][19] ), .op(
        n10498) );
  nor2_1 U12227 ( .ip1(n10494), .ip2(n10495), .op(n13427) );
  nand2_1 U12228 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][19] ), .op(
        n10497) );
  nor2_1 U12229 ( .ip1(n15315), .ip2(n10495), .op(n13428) );
  nand2_1 U12230 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][19] ), .op(
        n10496) );
  inv_1 U12231 ( .ip(\pipeline/imm[31] ), .op(n15324) );
  nor2_1 U12232 ( .ip1(n13209), .ip2(n10511), .op(n13445) );
  inv_1 U12233 ( .ip(n13445), .op(n10512) );
  or2_1 U12234 ( .ip1(n15324), .ip2(n10512), .op(n12503) );
  inv_1 U12235 ( .ip(n12503), .op(n12320) );
  inv_1 U12236 ( .ip(n17886), .op(n10513) );
  nand3_1 U12237 ( .ip1(\pipeline/inst_DX [2]), .ip2(n17786), .ip3(n10513), 
        .op(n12836) );
  nor2_1 U12238 ( .ip1(n15660), .ip2(n12836), .op(n10514) );
  nor2_1 U12239 ( .ip1(n12320), .ip2(n10514), .op(n10515) );
  nand2_1 U12240 ( .ip1(n10517), .ip2(n16552), .op(n10609) );
  nand2_1 U12241 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [18]), .op(n10520) );
  nand2_1 U12242 ( .ip1(\pipeline/alu_out_WB [18]), .ip2(n17895), .op(n10519)
         );
  nand2_1 U12243 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [18]), .op(
        n10518) );
  nand3_1 U12244 ( .ip1(n10520), .ip2(n10519), .ip3(n10518), .op(n18515) );
  nand2_1 U12245 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][18] ), .op(
        n10522) );
  nand2_1 U12246 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][18] ), .op(
        n10521) );
  nand2_1 U12247 ( .ip1(n10522), .ip2(n10521), .op(n10528) );
  nand2_1 U12248 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][18] ), .op(
        n10526) );
  nand2_1 U12249 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][18] ), .op(
        n10525) );
  nand2_1 U12250 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][18] ), .op(
        n10524) );
  nand2_1 U12251 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][18] ), .op(
        n10523) );
  not_ab_or_c_or_d U12252 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][18] ), .ip3(n10528), .ip4(n10527), .op(n10560) );
  nand2_1 U12253 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][18] ), .op(
        n10532) );
  nand2_1 U12254 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][18] ), .op(
        n10531) );
  nand2_1 U12255 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][18] ), .op(
        n10530) );
  nand2_1 U12256 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][18] ), .op(
        n10529) );
  and4_1 U12257 ( .ip1(n10532), .ip2(n10531), .ip3(n10530), .ip4(n10529), .op(
        n10559) );
  nand2_1 U12258 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][18] ), .op(
        n10536) );
  nand2_1 U12259 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][18] ), .op(
        n10535) );
  nand2_1 U12260 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][18] ), .op(
        n10534) );
  nand2_1 U12261 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][18] ), .op(
        n10533) );
  and4_1 U12262 ( .ip1(n10536), .ip2(n10535), .ip3(n10534), .ip4(n10533), .op(
        n10558) );
  nand2_1 U12263 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][18] ), .op(
        n10540) );
  nand2_1 U12264 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][18] ), .op(
        n10539) );
  nand2_1 U12265 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][18] ), .op(
        n10538) );
  nand2_1 U12266 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][18] ), .op(
        n10537) );
  nand2_1 U12267 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][18] ), .op(
        n10544) );
  nand2_1 U12268 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][18] ), .op(
        n10543) );
  nand2_1 U12269 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][18] ), .op(
        n10542) );
  nand2_1 U12270 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][18] ), .op(
        n10541) );
  nand2_1 U12271 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][18] ), .op(
        n10548) );
  nand2_1 U12272 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][18] ), .op(
        n10547) );
  nand2_1 U12273 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][18] ), .op(
        n10546) );
  nand2_1 U12274 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][18] ), .op(
        n10545) );
  nand2_1 U12275 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][18] ), .op(
        n10552) );
  nand2_1 U12276 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][18] ), .op(
        n10551) );
  nand2_1 U12277 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][18] ), .op(
        n10550) );
  nand2_1 U12278 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][18] ), .op(
        n10549) );
  mux2_1 U12279 ( .ip1(n18515), .ip2(n10561), .s(n10199), .op(n15597) );
  nand2_1 U12280 ( .ip1(n15597), .ip2(n13520), .op(n10563) );
  nand2_1 U12281 ( .ip1(n13521), .ip2(\pipeline/PC_DX [18]), .op(n10562) );
  nand2_2 U12282 ( .ip1(n10563), .ip2(n10562), .op(n16854) );
  nand2_1 U12283 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][18] ), .op(
        n10565) );
  nand2_1 U12284 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][18] ), .op(
        n10564) );
  nand2_1 U12285 ( .ip1(n10565), .ip2(n10564), .op(n10571) );
  nand2_1 U12286 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][18] ), .op(
        n10569) );
  nand2_1 U12287 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][18] ), .op(
        n10568) );
  nand2_1 U12288 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][18] ), .op(
        n10567) );
  nand2_1 U12289 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][18] ), .op(
        n10566) );
  not_ab_or_c_or_d U12290 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][18] ), .ip3(n10571), .ip4(n10570), .op(n10603) );
  nand2_1 U12291 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][18] ), .op(
        n10575) );
  nand2_1 U12292 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][18] ), .op(
        n10574) );
  nand2_1 U12293 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][18] ), .op(
        n10573) );
  nand2_1 U12294 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][18] ), .op(
        n10572) );
  and4_1 U12295 ( .ip1(n10575), .ip2(n10574), .ip3(n10573), .ip4(n10572), .op(
        n10602) );
  nand2_1 U12296 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][18] ), .op(
        n10579) );
  nand2_1 U12297 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][18] ), .op(
        n10578) );
  nand2_1 U12298 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][18] ), .op(
        n10577) );
  nand2_1 U12299 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][18] ), .op(
        n10576) );
  and4_1 U12300 ( .ip1(n10579), .ip2(n10578), .ip3(n10577), .ip4(n10576), .op(
        n10601) );
  nand2_1 U12301 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][18] ), .op(
        n10583) );
  nand2_1 U12302 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][18] ), .op(
        n10582) );
  nand2_1 U12303 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][18] ), .op(
        n10581) );
  nand2_1 U12304 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][18] ), .op(
        n10580) );
  nand2_1 U12305 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][18] ), .op(
        n10587) );
  nand2_1 U12306 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][18] ), .op(
        n10586) );
  nand2_1 U12307 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][18] ), .op(
        n10585) );
  nand2_1 U12308 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][18] ), .op(
        n10584) );
  nand2_1 U12309 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][18] ), .op(
        n10591) );
  nand2_1 U12310 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][18] ), .op(
        n10590) );
  nand2_1 U12311 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][18] ), .op(
        n10589) );
  nand2_1 U12312 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][18] ), .op(
        n10588) );
  nand2_1 U12313 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][18] ), .op(
        n10595) );
  nand2_1 U12314 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][18] ), .op(
        n10594) );
  nand2_1 U12315 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][18] ), .op(
        n10593) );
  nand2_1 U12316 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][18] ), .op(
        n10592) );
  nor2_1 U12317 ( .ip1(n15821), .ip2(n12836), .op(n10605) );
  nor2_1 U12318 ( .ip1(n12320), .ip2(n10605), .op(n10606) );
  nand2_1 U12319 ( .ip1(n10190), .ip2(n16557), .op(n13954) );
  nor2_1 U12320 ( .ip1(n13617), .ip2(n16552), .op(n10793) );
  or2_1 U12321 ( .ip1(n13954), .ip2(n10793), .op(n10608) );
  nand2_1 U12322 ( .ip1(n10609), .ip2(n10608), .op(n10610) );
  inv_1 U12323 ( .ip(n10610), .op(n10797) );
  nand2_1 U12324 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [17]), .op(n10613) );
  nand2_1 U12325 ( .ip1(\pipeline/alu_out_WB [17]), .ip2(n17895), .op(n10612)
         );
  nand2_1 U12326 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [17]), .op(
        n10611) );
  nand3_1 U12327 ( .ip1(n10613), .ip2(n10612), .ip3(n10611), .op(n19318) );
  nand2_1 U12328 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][17] ), .op(
        n10615) );
  nand2_1 U12329 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][17] ), .op(
        n10614) );
  nand2_1 U12330 ( .ip1(n10615), .ip2(n10614), .op(n10621) );
  nand2_1 U12331 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][17] ), .op(
        n10619) );
  nand2_1 U12332 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][17] ), .op(
        n10618) );
  nand2_1 U12333 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][17] ), .op(
        n10617) );
  nand2_1 U12334 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][17] ), .op(
        n10616) );
  not_ab_or_c_or_d U12335 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][17] ), .ip3(n10621), .ip4(n10620), .op(n10653) );
  nand2_1 U12336 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][17] ), .op(
        n10625) );
  nand2_1 U12337 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][17] ), .op(
        n10624) );
  nand2_1 U12338 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][17] ), .op(
        n10623) );
  nand2_1 U12339 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][17] ), .op(
        n10622) );
  and4_1 U12340 ( .ip1(n10625), .ip2(n10624), .ip3(n10623), .ip4(n10622), .op(
        n10652) );
  nand2_1 U12341 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][17] ), .op(
        n10629) );
  nand2_1 U12342 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][17] ), .op(
        n10628) );
  nand2_1 U12343 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][17] ), .op(
        n10627) );
  nand2_1 U12344 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][17] ), .op(
        n10626) );
  and4_1 U12345 ( .ip1(n10629), .ip2(n10628), .ip3(n10627), .ip4(n10626), .op(
        n10651) );
  nand2_1 U12346 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][17] ), .op(
        n10633) );
  nand2_1 U12347 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][17] ), .op(
        n10632) );
  nand2_1 U12348 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][17] ), .op(
        n10631) );
  nand2_1 U12349 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][17] ), .op(
        n10630) );
  nand2_1 U12350 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][17] ), .op(
        n10637) );
  nand2_1 U12351 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][17] ), .op(
        n10636) );
  nand2_1 U12352 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][17] ), .op(
        n10635) );
  nand2_1 U12353 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][17] ), .op(
        n10634) );
  nand2_1 U12354 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][17] ), .op(
        n10641) );
  nand2_1 U12355 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][17] ), .op(
        n10640) );
  nand2_1 U12356 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][17] ), .op(
        n10639) );
  nand2_1 U12357 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][17] ), .op(
        n10638) );
  nand2_1 U12358 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][17] ), .op(
        n10645) );
  nand2_1 U12359 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][17] ), .op(
        n10644) );
  nand2_1 U12360 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][17] ), .op(
        n10643) );
  nand2_1 U12361 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][17] ), .op(
        n10642) );
  mux2_1 U12362 ( .ip1(n19318), .ip2(n10654), .s(n10199), .op(n20007) );
  nand2_1 U12363 ( .ip1(n20007), .ip2(n13520), .op(n10656) );
  nand2_1 U12364 ( .ip1(n13521), .ip2(\pipeline/PC_DX [17]), .op(n10655) );
  nand2_1 U12365 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][17] ), .op(
        n10658) );
  nand2_1 U12366 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][17] ), .op(
        n10657) );
  nand2_1 U12367 ( .ip1(n10658), .ip2(n10657), .op(n10664) );
  nand2_1 U12368 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][17] ), .op(
        n10662) );
  nand2_1 U12369 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][17] ), .op(
        n10661) );
  nand2_1 U12370 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][17] ), .op(
        n10660) );
  nand2_1 U12371 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][17] ), .op(
        n10659) );
  not_ab_or_c_or_d U12372 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][17] ), .ip3(n10664), .ip4(n10663), .op(n10696) );
  nand2_1 U12373 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][17] ), .op(
        n10668) );
  nand2_1 U12374 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][17] ), .op(
        n10667) );
  nand2_1 U12375 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][17] ), .op(
        n10666) );
  nand2_1 U12376 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][17] ), .op(
        n10665) );
  and4_1 U12377 ( .ip1(n10668), .ip2(n10667), .ip3(n10666), .ip4(n10665), .op(
        n10695) );
  nand2_1 U12378 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][17] ), .op(
        n10672) );
  nand2_1 U12379 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][17] ), .op(
        n10671) );
  nand2_1 U12380 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][17] ), .op(
        n10670) );
  nand2_1 U12381 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][17] ), .op(
        n10669) );
  and4_1 U12382 ( .ip1(n10672), .ip2(n10671), .ip3(n10670), .ip4(n10669), .op(
        n10694) );
  nand2_1 U12383 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][17] ), .op(
        n10676) );
  nand2_1 U12384 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][17] ), .op(
        n10675) );
  nand2_1 U12385 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][17] ), .op(
        n10674) );
  nand2_1 U12386 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][17] ), .op(
        n10673) );
  nand2_1 U12387 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][17] ), .op(
        n10680) );
  nand2_1 U12388 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][17] ), .op(
        n10679) );
  nand2_1 U12389 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][17] ), .op(
        n10678) );
  nand2_1 U12390 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][17] ), .op(
        n10677) );
  nand2_1 U12391 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][17] ), .op(
        n10684) );
  nand2_1 U12392 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][17] ), .op(
        n10683) );
  nand2_1 U12393 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][17] ), .op(
        n10682) );
  nand2_1 U12394 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][17] ), .op(
        n10681) );
  nand2_1 U12395 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][17] ), .op(
        n10688) );
  nand2_1 U12396 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][17] ), .op(
        n10687) );
  nand2_1 U12397 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][17] ), .op(
        n10686) );
  nand2_1 U12398 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][17] ), .op(
        n10685) );
  mux2_1 U12399 ( .ip1(n19318), .ip2(n10697), .s(n12683), .op(n17387) );
  nor2_1 U12400 ( .ip1(n15782), .ip2(n12836), .op(n10698) );
  nor2_1 U12401 ( .ip1(n12320), .ip2(n10698), .op(n10699) );
  nand2_2 U12402 ( .ip1(n16627), .ip2(n16632), .op(n13885) );
  nand2_1 U12403 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [16]), .op(n10703) );
  nand2_1 U12404 ( .ip1(\pipeline/alu_out_WB [16]), .ip2(n17895), .op(n10702)
         );
  nand2_1 U12405 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [16]), .op(
        n10701) );
  nand3_1 U12406 ( .ip1(n10703), .ip2(n10702), .ip3(n10701), .op(n19323) );
  nand2_1 U12407 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][16] ), .op(
        n10705) );
  nand2_1 U12408 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][16] ), .op(
        n10704) );
  nand2_1 U12409 ( .ip1(n10705), .ip2(n10704), .op(n10711) );
  nand2_1 U12410 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][16] ), .op(
        n10709) );
  nand2_1 U12411 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][16] ), .op(
        n10708) );
  nand2_1 U12412 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][16] ), .op(
        n10707) );
  nand2_1 U12413 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][16] ), .op(
        n10706) );
  not_ab_or_c_or_d U12414 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][16] ), .ip3(n10711), .ip4(n10710), .op(n10743) );
  nand2_1 U12415 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][16] ), .op(
        n10715) );
  nand2_1 U12416 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][16] ), .op(
        n10714) );
  nand2_1 U12417 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][16] ), .op(
        n10713) );
  nand2_1 U12418 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][16] ), .op(
        n10712) );
  and4_1 U12419 ( .ip1(n10715), .ip2(n10714), .ip3(n10713), .ip4(n10712), .op(
        n10742) );
  nand2_1 U12420 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][16] ), .op(
        n10719) );
  nand2_1 U12421 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][16] ), .op(
        n10718) );
  nand2_1 U12422 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][16] ), .op(
        n10717) );
  nand2_1 U12423 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][16] ), .op(
        n10716) );
  and4_1 U12424 ( .ip1(n10719), .ip2(n10718), .ip3(n10717), .ip4(n10716), .op(
        n10741) );
  nand2_1 U12425 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][16] ), .op(
        n10723) );
  nand2_1 U12426 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][16] ), .op(
        n10722) );
  nand2_1 U12427 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][16] ), .op(
        n10721) );
  nand2_1 U12428 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][16] ), .op(
        n10720) );
  nand2_1 U12429 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][16] ), .op(
        n10727) );
  nand2_1 U12430 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][16] ), .op(
        n10726) );
  nand2_1 U12431 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][16] ), .op(
        n10725) );
  nand2_1 U12432 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][16] ), .op(
        n10724) );
  nand2_1 U12433 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][16] ), .op(
        n10731) );
  nand2_1 U12434 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][16] ), .op(
        n10730) );
  nand2_1 U12435 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][16] ), .op(
        n10729) );
  nand2_1 U12436 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][16] ), .op(
        n10728) );
  nand2_1 U12437 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][16] ), .op(
        n10735) );
  nand2_1 U12438 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][16] ), .op(
        n10734) );
  nand2_1 U12439 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][16] ), .op(
        n10733) );
  nand2_1 U12440 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][16] ), .op(
        n10732) );
  mux2_1 U12441 ( .ip1(n19323), .ip2(n10744), .s(n10199), .op(n14593) );
  nand2_1 U12442 ( .ip1(n14593), .ip2(n13520), .op(n10746) );
  nand2_1 U12443 ( .ip1(n13521), .ip2(\pipeline/PC_DX [16]), .op(n10745) );
  nor2_1 U12444 ( .ip1(n15833), .ip2(n12836), .op(n10747) );
  nor2_1 U12445 ( .ip1(n12320), .ip2(n10747), .op(n10790) );
  nand2_1 U12446 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][16] ), .op(
        n10749) );
  nand2_1 U12447 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][16] ), .op(
        n10748) );
  nand2_1 U12448 ( .ip1(n10749), .ip2(n10748), .op(n10755) );
  nand2_1 U12449 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][16] ), .op(
        n10753) );
  nand2_1 U12450 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][16] ), .op(
        n10752) );
  nand2_1 U12451 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][16] ), .op(
        n10751) );
  nand2_1 U12452 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][16] ), .op(
        n10750) );
  not_ab_or_c_or_d U12453 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][16] ), .ip3(n10755), .ip4(n10754), .op(n10787) );
  nand2_1 U12454 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][16] ), .op(
        n10759) );
  nand2_1 U12455 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][16] ), .op(
        n10758) );
  nand2_1 U12456 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][16] ), .op(
        n10757) );
  nand2_1 U12457 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][16] ), .op(
        n10756) );
  and4_1 U12458 ( .ip1(n10759), .ip2(n10758), .ip3(n10757), .ip4(n10756), .op(
        n10786) );
  nand2_1 U12459 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][16] ), .op(
        n10763) );
  nand2_1 U12460 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][16] ), .op(
        n10762) );
  nand2_1 U12461 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][16] ), .op(
        n10761) );
  nand2_1 U12462 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][16] ), .op(
        n10760) );
  and4_1 U12463 ( .ip1(n10763), .ip2(n10762), .ip3(n10761), .ip4(n10760), .op(
        n10785) );
  nand2_1 U12464 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][16] ), .op(
        n10767) );
  nand2_1 U12465 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][16] ), .op(
        n10766) );
  nand2_1 U12466 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][16] ), .op(
        n10765) );
  nand2_1 U12467 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][16] ), .op(
        n10764) );
  nand2_1 U12468 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][16] ), .op(
        n10771) );
  nand2_1 U12469 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][16] ), .op(
        n10770) );
  nand2_1 U12470 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][16] ), .op(
        n10769) );
  nand2_1 U12471 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][16] ), .op(
        n10768) );
  nand2_1 U12472 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][16] ), .op(
        n10775) );
  nand2_1 U12473 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][16] ), .op(
        n10774) );
  nand2_1 U12474 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][16] ), .op(
        n10773) );
  nand2_1 U12475 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][16] ), .op(
        n10772) );
  nand2_1 U12476 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][16] ), .op(
        n10779) );
  nand2_1 U12477 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][16] ), .op(
        n10778) );
  nand2_1 U12478 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][16] ), .op(
        n10777) );
  nand2_1 U12479 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][16] ), .op(
        n10776) );
  mux2_1 U12480 ( .ip1(n19323), .ip2(n10788), .s(n12683), .op(n22082) );
  nand2_1 U12481 ( .ip1(n22082), .ip2(n10201), .op(n10789) );
  inv_1 U12482 ( .ip(n16498), .op(n16418) );
  nand2_1 U12483 ( .ip1(n16526), .ip2(n16559), .op(n10791) );
  inv_1 U12484 ( .ip(n10190), .op(n16684) );
  nor2_1 U12485 ( .ip1(n10190), .ip2(n16557), .op(n10794) );
  nor2_1 U12486 ( .ip1(n10794), .ip2(n10793), .op(n13566) );
  nand2_1 U12487 ( .ip1(n10795), .ip2(n13566), .op(n10796) );
  nand2_1 U12488 ( .ip1(n10797), .ip2(n10796), .op(n13755) );
  nand2_1 U12489 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [22]), .op(n10800) );
  nand2_1 U12490 ( .ip1(\pipeline/alu_out_WB [22]), .ip2(n17895), .op(n10799)
         );
  nand2_1 U12491 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [22]), .op(
        n10798) );
  nand3_1 U12492 ( .ip1(n10800), .ip2(n10799), .ip3(n10798), .op(n19308) );
  buf_1 U12493 ( .ip(n11999), .op(n14057) );
  nand2_1 U12494 ( .ip1(n19308), .ip2(n12549), .op(n14059) );
  inv_1 U12495 ( .ip(n14059), .op(n10801) );
  nand2_1 U12496 ( .ip1(n13520), .ip2(n10801), .op(n10848) );
  nand2_1 U12497 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][22] ), .op(
        n10804) );
  nand2_1 U12498 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][22] ), .op(
        n10803) );
  nand2_1 U12499 ( .ip1(n10804), .ip2(n10803), .op(n10810) );
  nand2_1 U12500 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][22] ), .op(
        n10808) );
  nand2_1 U12501 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][22] ), .op(
        n10807) );
  nand2_1 U12502 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][22] ), .op(
        n10806) );
  nand2_1 U12503 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][22] ), .op(
        n10805) );
  not_ab_or_c_or_d U12504 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][22] ), .ip3(n10810), .ip4(n10809), .op(n10842) );
  nand2_1 U12505 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][22] ), .op(
        n10814) );
  nand2_1 U12506 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][22] ), .op(
        n10813) );
  nand2_1 U12507 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][22] ), .op(
        n10812) );
  nand2_1 U12508 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][22] ), .op(
        n10811) );
  and4_1 U12509 ( .ip1(n10814), .ip2(n10813), .ip3(n10812), .ip4(n10811), .op(
        n10841) );
  nand2_1 U12510 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][22] ), .op(
        n10818) );
  nand2_1 U12511 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][22] ), .op(
        n10817) );
  nand2_1 U12512 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][22] ), .op(
        n10816) );
  nand2_1 U12513 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][22] ), .op(
        n10815) );
  and4_1 U12514 ( .ip1(n10818), .ip2(n10817), .ip3(n10816), .ip4(n10815), .op(
        n10840) );
  nand2_1 U12515 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][22] ), .op(
        n10822) );
  nand2_1 U12516 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][22] ), .op(
        n10821) );
  nand2_1 U12517 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][22] ), .op(
        n10820) );
  nand2_1 U12518 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][22] ), .op(
        n10819) );
  nand2_1 U12519 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][22] ), .op(
        n10826) );
  nand2_1 U12520 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][22] ), .op(
        n10825) );
  nand2_1 U12521 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][22] ), .op(
        n10824) );
  nand2_1 U12522 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][22] ), .op(
        n10823) );
  nand2_1 U12523 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][22] ), .op(
        n10830) );
  nand2_1 U12524 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][22] ), .op(
        n10829) );
  nand2_1 U12525 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][22] ), .op(
        n10828) );
  nand2_1 U12526 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][22] ), .op(
        n10827) );
  nand2_1 U12527 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][22] ), .op(
        n10834) );
  nand2_1 U12528 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][22] ), .op(
        n10833) );
  nand2_1 U12529 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][22] ), .op(
        n10832) );
  nand2_1 U12530 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][22] ), .op(
        n10831) );
  inv_1 U12531 ( .ip(n14056), .op(n10843) );
  nor2_1 U12532 ( .ip1(n10511), .ip2(n10843), .op(n10844) );
  nand2_1 U12533 ( .ip1(n13162), .ip2(n10844), .op(n10845) );
  inv_1 U12534 ( .ip(n10845), .op(n10846) );
  nor2_1 U12535 ( .ip1(n10802), .ip2(n10846), .op(n10847) );
  nand2_1 U12536 ( .ip1(n10201), .ip2(n19308), .op(n10850) );
  inv_1 U12537 ( .ip(n10850), .op(n10851) );
  nand2_1 U12538 ( .ip1(n12880), .ip2(n10851), .op(n10897) );
  nand2_1 U12539 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][22] ), .op(
        n10853) );
  nand2_1 U12540 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][22] ), .op(
        n10852) );
  nand2_1 U12541 ( .ip1(n10853), .ip2(n10852), .op(n10859) );
  nand2_1 U12542 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][22] ), .op(
        n10857) );
  nand2_1 U12543 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][22] ), .op(
        n10856) );
  nand2_1 U12544 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][22] ), .op(
        n10855) );
  nand2_1 U12545 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][22] ), .op(
        n10854) );
  not_ab_or_c_or_d U12546 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][22] ), .ip3(n10859), .ip4(n10858), .op(n10891) );
  nand2_1 U12547 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][22] ), .op(
        n10863) );
  nand2_1 U12548 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][22] ), .op(
        n10862) );
  nand2_1 U12549 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][22] ), .op(
        n10861) );
  nand2_1 U12550 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][22] ), .op(
        n10860) );
  and4_1 U12551 ( .ip1(n10863), .ip2(n10862), .ip3(n10861), .ip4(n10860), .op(
        n10890) );
  nand2_1 U12552 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][22] ), .op(
        n10867) );
  nand2_1 U12553 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][22] ), .op(
        n10866) );
  nand2_1 U12554 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][22] ), .op(
        n10865) );
  nand2_1 U12555 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][22] ), .op(
        n10864) );
  and4_1 U12556 ( .ip1(n10867), .ip2(n10866), .ip3(n10865), .ip4(n10864), .op(
        n10889) );
  nand2_1 U12557 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][22] ), .op(
        n10871) );
  nand2_1 U12558 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][22] ), .op(
        n10870) );
  nand2_1 U12559 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][22] ), .op(
        n10869) );
  nand2_1 U12560 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][22] ), .op(
        n10868) );
  nand2_1 U12561 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][22] ), .op(
        n10875) );
  nand2_1 U12562 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][22] ), .op(
        n10874) );
  nand2_1 U12563 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][22] ), .op(
        n10873) );
  nand2_1 U12564 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][22] ), .op(
        n10872) );
  nand2_1 U12565 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][22] ), .op(
        n10879) );
  nand2_1 U12566 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][22] ), .op(
        n10878) );
  nand2_1 U12567 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][22] ), .op(
        n10877) );
  nand2_1 U12568 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][22] ), .op(
        n10876) );
  nand2_1 U12569 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][22] ), .op(
        n10883) );
  nand2_1 U12570 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][22] ), .op(
        n10882) );
  nand2_1 U12571 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][22] ), .op(
        n10881) );
  nand2_1 U12572 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][22] ), .op(
        n10880) );
  and2_1 U12573 ( .ip1(n17398), .ip2(n10201), .op(n10892) );
  nand2_1 U12574 ( .ip1(n13315), .ip2(n10892), .op(n10895) );
  inv_1 U12575 ( .ip(\pipeline/inst_DX [22]), .op(n13207) );
  nor2_1 U12576 ( .ip1(n13207), .ip2(n12836), .op(n10893) );
  nor2_1 U12577 ( .ip1(n12320), .ip2(n10893), .op(n10894) );
  nand2_1 U12578 ( .ip1(n10897), .ip2(n10896), .op(n17173) );
  nor2_1 U12579 ( .ip1(n10849), .ip2(n17173), .op(n10991) );
  nand2_1 U12580 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [23]), .op(n10900) );
  nand2_1 U12581 ( .ip1(\pipeline/alu_out_WB [23]), .ip2(n17895), .op(n10899)
         );
  nand2_1 U12582 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [23]), .op(
        n10898) );
  nand3_1 U12583 ( .ip1(n10900), .ip2(n10899), .ip3(n10898), .op(n19301) );
  nand2_1 U12584 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][23] ), .op(
        n10902) );
  nand2_1 U12585 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][23] ), .op(
        n10901) );
  nand2_1 U12586 ( .ip1(n10902), .ip2(n10901), .op(n10908) );
  nand2_1 U12587 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][23] ), .op(
        n10906) );
  nand2_1 U12588 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][23] ), .op(
        n10905) );
  nand2_1 U12589 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][23] ), .op(
        n10904) );
  nand2_1 U12590 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][23] ), .op(
        n10903) );
  not_ab_or_c_or_d U12591 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][23] ), .ip3(n10908), .ip4(n10907), .op(n10940) );
  nand2_1 U12592 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][23] ), .op(
        n10912) );
  nand2_1 U12593 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][23] ), .op(
        n10911) );
  nand2_1 U12594 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][23] ), .op(
        n10910) );
  nand2_1 U12595 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][23] ), .op(
        n10909) );
  and4_1 U12596 ( .ip1(n10912), .ip2(n10911), .ip3(n10910), .ip4(n10909), .op(
        n10939) );
  nand2_1 U12597 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][23] ), .op(
        n10916) );
  nand2_1 U12598 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][23] ), .op(
        n10915) );
  nand2_1 U12599 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][23] ), .op(
        n10914) );
  nand2_1 U12600 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][23] ), .op(
        n10913) );
  and4_1 U12601 ( .ip1(n10916), .ip2(n10915), .ip3(n10914), .ip4(n10913), .op(
        n10938) );
  nand2_1 U12602 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][23] ), .op(
        n10920) );
  nand2_1 U12603 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][23] ), .op(
        n10919) );
  nand2_1 U12604 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][23] ), .op(
        n10918) );
  nand2_1 U12605 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][23] ), .op(
        n10917) );
  nand2_1 U12606 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][23] ), .op(
        n10924) );
  nand2_1 U12607 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][23] ), .op(
        n10923) );
  nand2_1 U12608 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][23] ), .op(
        n10922) );
  nand2_1 U12609 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][23] ), .op(
        n10921) );
  nand2_1 U12610 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][23] ), .op(
        n10928) );
  nand2_1 U12611 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][23] ), .op(
        n10927) );
  nand2_1 U12612 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][23] ), .op(
        n10926) );
  nand2_1 U12613 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][23] ), .op(
        n10925) );
  nand2_1 U12614 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][23] ), .op(
        n10932) );
  nand2_1 U12615 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][23] ), .op(
        n10931) );
  nand2_1 U12616 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][23] ), .op(
        n10930) );
  nand2_1 U12617 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][23] ), .op(
        n10929) );
  mux2_1 U12618 ( .ip1(n19301), .ip2(n10941), .s(n10199), .op(n15401) );
  nand2_1 U12619 ( .ip1(n15401), .ip2(n13520), .op(n10943) );
  nand2_1 U12620 ( .ip1(n13521), .ip2(\pipeline/PC_DX [23]), .op(n10942) );
  inv_1 U12621 ( .ip(n13654), .op(n18738) );
  nand2_1 U12622 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][23] ), .op(
        n10946) );
  nand2_1 U12623 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][23] ), .op(
        n10945) );
  nand2_1 U12624 ( .ip1(n10946), .ip2(n10945), .op(n10952) );
  nand2_1 U12625 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][23] ), .op(
        n10950) );
  nand2_1 U12626 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][23] ), .op(
        n10949) );
  nand2_1 U12627 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][23] ), .op(
        n10948) );
  nand2_1 U12628 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][23] ), .op(
        n10947) );
  not_ab_or_c_or_d U12629 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][23] ), .ip3(n10952), .ip4(n10951), .op(n10984) );
  nand2_1 U12630 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][23] ), .op(
        n10956) );
  nand2_1 U12631 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][23] ), .op(
        n10955) );
  nand2_1 U12632 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][23] ), .op(
        n10954) );
  nand2_1 U12633 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][23] ), .op(
        n10953) );
  and4_1 U12634 ( .ip1(n10956), .ip2(n10955), .ip3(n10954), .ip4(n10953), .op(
        n10983) );
  nand2_1 U12635 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][23] ), .op(
        n10960) );
  nand2_1 U12636 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][23] ), .op(
        n10959) );
  nand2_1 U12637 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][23] ), .op(
        n10958) );
  nand2_1 U12638 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][23] ), .op(
        n10957) );
  and4_1 U12639 ( .ip1(n10960), .ip2(n10959), .ip3(n10958), .ip4(n10957), .op(
        n10982) );
  nand2_1 U12640 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][23] ), .op(
        n10964) );
  nand2_1 U12641 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][23] ), .op(
        n10963) );
  nand2_1 U12642 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][23] ), .op(
        n10962) );
  nand2_1 U12643 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][23] ), .op(
        n10961) );
  nand2_1 U12644 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][23] ), .op(
        n10968) );
  nand2_1 U12645 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][23] ), .op(
        n10967) );
  nand2_1 U12646 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][23] ), .op(
        n10966) );
  nand2_1 U12647 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][23] ), .op(
        n10965) );
  nand2_1 U12648 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][23] ), .op(
        n10972) );
  nand2_1 U12649 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][23] ), .op(
        n10971) );
  nand2_1 U12650 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][23] ), .op(
        n10970) );
  nand2_1 U12651 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][23] ), .op(
        n10969) );
  nand2_1 U12652 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][23] ), .op(
        n10976) );
  nand2_1 U12653 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][23] ), .op(
        n10975) );
  nand2_1 U12654 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][23] ), .op(
        n10974) );
  nand2_1 U12655 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][23] ), .op(
        n10973) );
  and4_1 U12656 ( .ip1(n10984), .ip2(n10983), .ip3(n10982), .ip4(n10981), .op(
        n10985) );
  or2_1 U12657 ( .ip1(n13315), .ip2(n19301), .op(n17405) );
  nand2_1 U12658 ( .ip1(n17405), .ip2(n10201), .op(n10986) );
  inv_1 U12659 ( .ip(n10986), .op(n10987) );
  nor2_1 U12660 ( .ip1(n13117), .ip2(n12836), .op(n10988) );
  nor2_1 U12661 ( .ip1(n12320), .ip2(n10988), .op(n10989) );
  nor2_1 U12662 ( .ip1(n13654), .ip2(n16594), .op(n11176) );
  nor2_1 U12663 ( .ip1(n10991), .ip2(n11176), .op(n11184) );
  nand2_1 U12664 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][20] ), .op(
        n10993) );
  nand2_1 U12665 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][20] ), .op(
        n10992) );
  nand2_1 U12666 ( .ip1(n10993), .ip2(n10992), .op(n10999) );
  nand2_1 U12667 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][20] ), .op(
        n10997) );
  nand2_1 U12668 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][20] ), .op(
        n10996) );
  nand2_1 U12669 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][20] ), .op(
        n10995) );
  nand2_1 U12670 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][20] ), .op(
        n10994) );
  not_ab_or_c_or_d U12671 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][20] ), .ip3(n10999), .ip4(n10998), .op(n11031) );
  nand2_1 U12672 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][20] ), .op(
        n11003) );
  nand2_1 U12673 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][20] ), .op(
        n11002) );
  nand2_1 U12674 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][20] ), .op(
        n11001) );
  nand2_1 U12675 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][20] ), .op(
        n11000) );
  and4_1 U12676 ( .ip1(n11003), .ip2(n11002), .ip3(n11001), .ip4(n11000), .op(
        n11030) );
  nand2_1 U12677 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][20] ), .op(
        n11007) );
  nand2_1 U12678 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][20] ), .op(
        n11006) );
  nand2_1 U12679 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][20] ), .op(
        n11005) );
  nand2_1 U12680 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][20] ), .op(
        n11004) );
  and4_1 U12681 ( .ip1(n11007), .ip2(n11006), .ip3(n11005), .ip4(n11004), .op(
        n11029) );
  nand2_1 U12682 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][20] ), .op(
        n11011) );
  nand2_1 U12683 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][20] ), .op(
        n11010) );
  nand2_1 U12684 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][20] ), .op(
        n11009) );
  nand2_1 U12685 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][20] ), .op(
        n11008) );
  nand2_1 U12686 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][20] ), .op(
        n11015) );
  nand2_1 U12687 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][20] ), .op(
        n11014) );
  nand2_1 U12688 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][20] ), .op(
        n11013) );
  nand2_1 U12689 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][20] ), .op(
        n11012) );
  nand2_1 U12690 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][20] ), .op(
        n11019) );
  nand2_1 U12691 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][20] ), .op(
        n11018) );
  nand2_1 U12692 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][20] ), .op(
        n11017) );
  nand2_1 U12693 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][20] ), .op(
        n11016) );
  nand2_1 U12694 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][20] ), .op(
        n11023) );
  nand2_1 U12695 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][20] ), .op(
        n11022) );
  nand2_1 U12696 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][20] ), .op(
        n11021) );
  nand2_1 U12697 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][20] ), .op(
        n11020) );
  nand2_1 U12698 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [20]), .op(n11034) );
  nand2_1 U12699 ( .ip1(\pipeline/alu_out_WB [20]), .ip2(n17895), .op(n11033)
         );
  nand2_1 U12700 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [20]), .op(
        n11032) );
  nand3_1 U12701 ( .ip1(n11034), .ip2(n11033), .ip3(n11032), .op(n19313) );
  inv_1 U12702 ( .ip(n13364), .op(n12549) );
  mux2_1 U12703 ( .ip1(n11035), .ip2(n19313), .s(n12549), .op(n15356) );
  nand2_1 U12704 ( .ip1(n15356), .ip2(n13520), .op(n11037) );
  nand2_1 U12705 ( .ip1(n13521), .ip2(\pipeline/PC_DX [20]), .op(n11036) );
  nand2_1 U12706 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][20] ), .op(
        n11039) );
  nand2_1 U12707 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][20] ), .op(
        n11038) );
  nand2_1 U12708 ( .ip1(n11039), .ip2(n11038), .op(n11045) );
  nand2_1 U12709 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][20] ), .op(
        n11043) );
  nand2_1 U12710 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][20] ), .op(
        n11042) );
  nand2_1 U12711 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][20] ), .op(
        n11041) );
  nand2_1 U12712 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][20] ), .op(
        n11040) );
  not_ab_or_c_or_d U12713 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][20] ), .ip3(n11045), .ip4(n11044), .op(n11077) );
  nand2_1 U12714 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][20] ), .op(
        n11049) );
  nand2_1 U12715 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][20] ), .op(
        n11048) );
  nand2_1 U12716 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][20] ), .op(
        n11047) );
  nand2_1 U12717 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][20] ), .op(
        n11046) );
  and4_1 U12718 ( .ip1(n11049), .ip2(n11048), .ip3(n11047), .ip4(n11046), .op(
        n11076) );
  nand2_1 U12719 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][20] ), .op(
        n11053) );
  nand2_1 U12720 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][20] ), .op(
        n11052) );
  nand2_1 U12721 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][20] ), .op(
        n11051) );
  nand2_1 U12722 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][20] ), .op(
        n11050) );
  and4_1 U12723 ( .ip1(n11053), .ip2(n11052), .ip3(n11051), .ip4(n11050), .op(
        n11075) );
  nand2_1 U12724 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][20] ), .op(
        n11057) );
  nand2_1 U12725 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][20] ), .op(
        n11056) );
  nand2_1 U12726 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][20] ), .op(
        n11055) );
  nand2_1 U12727 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][20] ), .op(
        n11054) );
  nand2_1 U12728 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][20] ), .op(
        n11061) );
  nand2_1 U12729 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][20] ), .op(
        n11060) );
  nand2_1 U12730 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][20] ), .op(
        n11059) );
  nand2_1 U12731 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][20] ), .op(
        n11058) );
  nand2_1 U12732 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][20] ), .op(
        n11065) );
  nand2_1 U12733 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][20] ), .op(
        n11064) );
  nand2_1 U12734 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][20] ), .op(
        n11063) );
  nand2_1 U12735 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][20] ), .op(
        n11062) );
  nand2_1 U12736 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][20] ), .op(
        n11069) );
  nand2_1 U12737 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][20] ), .op(
        n11068) );
  nand2_1 U12738 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][20] ), .op(
        n11067) );
  nand2_1 U12739 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][20] ), .op(
        n11066) );
  mux2_1 U12740 ( .ip1(n19313), .ip2(n11078), .s(n13441), .op(n22085) );
  nand2_1 U12741 ( .ip1(n22085), .ip2(n10201), .op(n11082) );
  nor2_1 U12742 ( .ip1(n11079), .ip2(n12836), .op(n11080) );
  nor2_1 U12743 ( .ip1(n12320), .ip2(n11080), .op(n11081) );
  nand2_1 U12744 ( .ip1(n11082), .ip2(n11081), .op(n16550) );
  nor2_1 U12745 ( .ip1(n11180), .ip2(n16550), .op(n11173) );
  nand2_1 U12746 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [21]), .op(n11085) );
  nand2_1 U12747 ( .ip1(\pipeline/alu_out_WB [21]), .ip2(n17895), .op(n11084)
         );
  nand2_1 U12748 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [21]), .op(
        n11083) );
  nand3_1 U12749 ( .ip1(n11085), .ip2(n11084), .ip3(n11083), .op(n18646) );
  nand2_1 U12750 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][21] ), .op(
        n11087) );
  nand2_1 U12751 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][21] ), .op(
        n11086) );
  nand2_1 U12752 ( .ip1(n11087), .ip2(n11086), .op(n11093) );
  nand2_1 U12753 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][21] ), .op(
        n11091) );
  nand2_1 U12754 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][21] ), .op(
        n11090) );
  nand2_1 U12755 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][21] ), .op(
        n11089) );
  nand2_1 U12756 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][21] ), .op(
        n11088) );
  not_ab_or_c_or_d U12757 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][21] ), .ip3(n11093), .ip4(n11092), .op(n11125) );
  nand2_1 U12758 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][21] ), .op(
        n11097) );
  nand2_1 U12759 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][21] ), .op(
        n11096) );
  nand2_1 U12760 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][21] ), .op(
        n11095) );
  nand2_1 U12761 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][21] ), .op(
        n11094) );
  and4_1 U12762 ( .ip1(n11097), .ip2(n11096), .ip3(n11095), .ip4(n11094), .op(
        n11124) );
  nand2_1 U12763 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][21] ), .op(
        n11101) );
  nand2_1 U12764 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][21] ), .op(
        n11100) );
  nand2_1 U12765 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][21] ), .op(
        n11099) );
  nand2_1 U12766 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][21] ), .op(
        n11098) );
  and4_1 U12767 ( .ip1(n11101), .ip2(n11100), .ip3(n11099), .ip4(n11098), .op(
        n11123) );
  nand2_1 U12768 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][21] ), .op(
        n11105) );
  nand2_1 U12769 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][21] ), .op(
        n11104) );
  nand2_1 U12770 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][21] ), .op(
        n11103) );
  nand2_1 U12771 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][21] ), .op(
        n11102) );
  nand2_1 U12772 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][21] ), .op(
        n11109) );
  nand2_1 U12773 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][21] ), .op(
        n11108) );
  nand2_1 U12774 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][21] ), .op(
        n11107) );
  nand2_1 U12775 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][21] ), .op(
        n11106) );
  nand2_1 U12776 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][21] ), .op(
        n11113) );
  nand2_1 U12777 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][21] ), .op(
        n11112) );
  nand2_1 U12778 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][21] ), .op(
        n11111) );
  nand2_1 U12779 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][21] ), .op(
        n11110) );
  nand2_1 U12780 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][21] ), .op(
        n11117) );
  nand2_1 U12781 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][21] ), .op(
        n11116) );
  nand2_1 U12782 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][21] ), .op(
        n11115) );
  nand2_1 U12783 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][21] ), .op(
        n11114) );
  mux2_1 U12784 ( .ip1(n18646), .ip2(n11126), .s(n10199), .op(n20586) );
  nand2_1 U12785 ( .ip1(n20586), .ip2(n13520), .op(n11128) );
  nand2_1 U12786 ( .ip1(n13521), .ip2(\pipeline/PC_DX [21]), .op(n11127) );
  or2_1 U12787 ( .ip1(n13315), .ip2(n18646), .op(n17392) );
  nand2_1 U12788 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][21] ), .op(
        n11130) );
  nand2_1 U12789 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][21] ), .op(
        n11129) );
  nand2_1 U12790 ( .ip1(n11130), .ip2(n11129), .op(n11136) );
  nand2_1 U12791 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][21] ), .op(
        n11134) );
  nand2_1 U12792 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][21] ), .op(
        n11133) );
  nand2_1 U12793 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][21] ), .op(
        n11132) );
  nand2_1 U12794 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][21] ), .op(
        n11131) );
  not_ab_or_c_or_d U12795 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][21] ), .ip3(n11136), .ip4(n11135), .op(n11168) );
  nand2_1 U12796 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][21] ), .op(
        n11140) );
  nand2_1 U12797 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][21] ), .op(
        n11139) );
  nand2_1 U12798 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][21] ), .op(
        n11138) );
  nand2_1 U12799 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][21] ), .op(
        n11137) );
  and4_1 U12800 ( .ip1(n11140), .ip2(n11139), .ip3(n11138), .ip4(n11137), .op(
        n11167) );
  nand2_1 U12801 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][21] ), .op(
        n11144) );
  nand2_1 U12802 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][21] ), .op(
        n11143) );
  nand2_1 U12803 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][21] ), .op(
        n11142) );
  nand2_1 U12804 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][21] ), .op(
        n11141) );
  and4_1 U12805 ( .ip1(n11144), .ip2(n11143), .ip3(n11142), .ip4(n11141), .op(
        n11166) );
  nand2_1 U12806 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][21] ), .op(
        n11148) );
  nand2_1 U12807 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][21] ), .op(
        n11147) );
  nand2_1 U12808 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][21] ), .op(
        n11146) );
  nand2_1 U12809 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][21] ), .op(
        n11145) );
  nand2_1 U12810 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][21] ), .op(
        n11152) );
  nand2_1 U12811 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][21] ), .op(
        n11151) );
  nand2_1 U12812 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][21] ), .op(
        n11150) );
  nand2_1 U12813 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][21] ), .op(
        n11149) );
  nand2_1 U12814 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][21] ), .op(
        n11156) );
  nand2_1 U12815 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][21] ), .op(
        n11155) );
  nand2_1 U12816 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][21] ), .op(
        n11154) );
  nand2_1 U12817 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][21] ), .op(
        n11153) );
  nand2_1 U12818 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][21] ), .op(
        n11160) );
  nand2_1 U12819 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][21] ), .op(
        n11159) );
  nand2_1 U12820 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][21] ), .op(
        n11158) );
  nand2_1 U12821 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][21] ), .op(
        n11157) );
  and4_1 U12822 ( .ip1(n11168), .ip2(n11167), .ip3(n11166), .ip4(n11165), .op(
        n11169) );
  nand2_1 U12823 ( .ip1(n11169), .ip2(n13315), .op(n17391) );
  nand3_1 U12824 ( .ip1(n17392), .ip2(n10201), .ip3(n17391), .op(n11172) );
  nor2_1 U12825 ( .ip1(n13319), .ip2(n12836), .op(n11170) );
  nor2_1 U12826 ( .ip1(n12320), .ip2(n11170), .op(n11171) );
  nand2_1 U12827 ( .ip1(n11172), .ip2(n11171), .op(n16545) );
  nor2_1 U12828 ( .ip1(n10192), .ip2(n16545), .op(n11181) );
  nor2_1 U12829 ( .ip1(n11173), .ip2(n11181), .op(n11174) );
  nand2_1 U12830 ( .ip1(n11184), .ip2(n11174), .op(n13569) );
  inv_1 U12831 ( .ip(n13569), .op(n11175) );
  nand2_1 U12832 ( .ip1(n13755), .ip2(n11175), .op(n11189) );
  nand2_1 U12833 ( .ip1(n13654), .ip2(n16594), .op(n11179) );
  nand2_1 U12834 ( .ip1(n10849), .ip2(n17173), .op(n11177) );
  or2_1 U12835 ( .ip1(n11177), .ip2(n11176), .op(n11178) );
  nand2_1 U12836 ( .ip1(n11179), .ip2(n11178), .op(n11187) );
  nand2_1 U12837 ( .ip1(n10192), .ip2(n16545), .op(n11183) );
  nand2_1 U12838 ( .ip1(n11180), .ip2(n16550), .op(n13906) );
  or2_1 U12839 ( .ip1(n13906), .ip2(n11181), .op(n11182) );
  nand2_1 U12840 ( .ip1(n11183), .ip2(n11182), .op(n11185) );
  and2_1 U12841 ( .ip1(n11185), .ip2(n11184), .op(n11186) );
  nor2_1 U12842 ( .ip1(n11187), .ip2(n11186), .op(n11188) );
  nand2_1 U12843 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [27]), .op(n11192) );
  nand2_1 U12844 ( .ip1(\pipeline/alu_out_WB [27]), .ip2(n17895), .op(n11191)
         );
  nand2_1 U12845 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [27]), .op(
        n11190) );
  nand3_1 U12846 ( .ip1(n11192), .ip2(n11191), .ip3(n11190), .op(n19166) );
  nand2_1 U12847 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][27] ), .op(
        n11194) );
  nand2_1 U12848 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][27] ), .op(
        n11193) );
  nand2_1 U12849 ( .ip1(n11194), .ip2(n11193), .op(n11200) );
  nand2_1 U12850 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][27] ), .op(
        n11198) );
  nand2_1 U12851 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][27] ), .op(
        n11197) );
  nand2_1 U12852 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][27] ), .op(
        n11196) );
  nand2_1 U12853 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][27] ), .op(
        n11195) );
  not_ab_or_c_or_d U12854 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][27] ), .ip3(n11200), .ip4(n11199), .op(n11232) );
  nand2_1 U12855 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][27] ), .op(
        n11204) );
  nand2_1 U12856 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][27] ), .op(
        n11203) );
  nand2_1 U12857 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][27] ), .op(
        n11202) );
  nand2_1 U12858 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][27] ), .op(
        n11201) );
  and4_1 U12859 ( .ip1(n11204), .ip2(n11203), .ip3(n11202), .ip4(n11201), .op(
        n11231) );
  nand2_1 U12860 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][27] ), .op(
        n11208) );
  nand2_1 U12861 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][27] ), .op(
        n11207) );
  nand2_1 U12862 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][27] ), .op(
        n11206) );
  nand2_1 U12863 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][27] ), .op(
        n11205) );
  and4_1 U12864 ( .ip1(n11208), .ip2(n11207), .ip3(n11206), .ip4(n11205), .op(
        n11230) );
  nand2_1 U12865 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][27] ), .op(
        n11212) );
  nand2_1 U12866 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][27] ), .op(
        n11211) );
  nand2_1 U12867 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][27] ), .op(
        n11210) );
  nand2_1 U12868 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][27] ), .op(
        n11209) );
  nand2_1 U12869 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][27] ), .op(
        n11216) );
  nand2_1 U12870 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][27] ), .op(
        n11215) );
  nand2_1 U12871 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][27] ), .op(
        n11214) );
  nand2_1 U12872 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][27] ), .op(
        n11213) );
  nand2_1 U12873 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][27] ), .op(
        n11220) );
  nand2_1 U12874 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][27] ), .op(
        n11219) );
  nand2_1 U12875 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][27] ), .op(
        n11218) );
  nand2_1 U12876 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][27] ), .op(
        n11217) );
  nand2_1 U12877 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][27] ), .op(
        n11224) );
  nand2_1 U12878 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][27] ), .op(
        n11223) );
  nand2_1 U12879 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][27] ), .op(
        n11222) );
  nand2_1 U12880 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][27] ), .op(
        n11221) );
  mux2_1 U12881 ( .ip1(n19166), .ip2(n11233), .s(n10200), .op(n16237) );
  nand2_1 U12882 ( .ip1(n16237), .ip2(n13520), .op(n11235) );
  nand2_1 U12883 ( .ip1(n13521), .ip2(\pipeline/PC_DX [27]), .op(n11234) );
  nand2_1 U12884 ( .ip1(n11235), .ip2(n11234), .op(n13742) );
  nand2_1 U12885 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][27] ), .op(
        n11237) );
  nand2_1 U12886 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][27] ), .op(
        n11236) );
  nand2_1 U12887 ( .ip1(n11237), .ip2(n11236), .op(n11243) );
  nand2_1 U12888 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][27] ), .op(
        n11241) );
  nand2_1 U12889 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][27] ), .op(
        n11240) );
  nand2_1 U12890 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][27] ), .op(
        n11239) );
  nand2_1 U12891 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][27] ), .op(
        n11238) );
  not_ab_or_c_or_d U12892 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][27] ), .ip3(n11243), .ip4(n11242), .op(n11275) );
  nand2_1 U12893 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][27] ), .op(
        n11247) );
  nand2_1 U12894 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][27] ), .op(
        n11246) );
  nand2_1 U12895 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][27] ), .op(
        n11245) );
  nand2_1 U12896 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][27] ), .op(
        n11244) );
  and4_1 U12897 ( .ip1(n11247), .ip2(n11246), .ip3(n11245), .ip4(n11244), .op(
        n11274) );
  nand2_1 U12898 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][27] ), .op(
        n11251) );
  nand2_1 U12899 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][27] ), .op(
        n11250) );
  nand2_1 U12900 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][27] ), .op(
        n11249) );
  nand2_1 U12901 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][27] ), .op(
        n11248) );
  and4_1 U12902 ( .ip1(n11251), .ip2(n11250), .ip3(n11249), .ip4(n11248), .op(
        n11273) );
  nand2_1 U12903 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][27] ), .op(
        n11255) );
  nand2_1 U12904 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][27] ), .op(
        n11254) );
  nand2_1 U12905 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][27] ), .op(
        n11253) );
  nand2_1 U12906 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][27] ), .op(
        n11252) );
  nand2_1 U12907 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][27] ), .op(
        n11259) );
  nand2_1 U12908 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][27] ), .op(
        n11258) );
  nand2_1 U12909 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][27] ), .op(
        n11257) );
  nand2_1 U12910 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][27] ), .op(
        n11256) );
  nand2_1 U12911 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][27] ), .op(
        n11263) );
  nand2_1 U12912 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][27] ), .op(
        n11262) );
  nand2_1 U12913 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][27] ), .op(
        n11261) );
  nand2_1 U12914 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][27] ), .op(
        n11260) );
  nand2_1 U12915 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][27] ), .op(
        n11267) );
  nand2_1 U12916 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][27] ), .op(
        n11266) );
  nand2_1 U12917 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][27] ), .op(
        n11265) );
  nand2_1 U12918 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][27] ), .op(
        n11264) );
  mux2_1 U12919 ( .ip1(n19166), .ip2(n11276), .s(n12683), .op(n21277) );
  nand2_1 U12920 ( .ip1(n21277), .ip2(n10201), .op(n11279) );
  nor2_1 U12921 ( .ip1(n15339), .ip2(n12836), .op(n11277) );
  nor2_1 U12922 ( .ip1(n12320), .ip2(n11277), .op(n11278) );
  inv_1 U12923 ( .ip(n13601), .op(n13743) );
  nand2_1 U12924 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [26]), .op(n11282) );
  nand2_1 U12925 ( .ip1(\pipeline/alu_out_WB [26]), .ip2(n17895), .op(n11281)
         );
  nand2_1 U12926 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [26]), .op(
        n11280) );
  nand3_1 U12927 ( .ip1(n11282), .ip2(n11281), .ip3(n11280), .op(n19089) );
  nand2_1 U12928 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][26] ), .op(
        n11284) );
  nand2_1 U12929 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][26] ), .op(
        n11283) );
  nand2_1 U12930 ( .ip1(n11284), .ip2(n11283), .op(n11290) );
  nand2_1 U12931 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][26] ), .op(
        n11288) );
  nand2_1 U12932 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][26] ), .op(
        n11287) );
  nand2_1 U12933 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][26] ), .op(
        n11286) );
  nand2_1 U12934 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][26] ), .op(
        n11285) );
  not_ab_or_c_or_d U12935 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][26] ), .ip3(n11290), .ip4(n11289), .op(n11322) );
  nand2_1 U12936 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][26] ), .op(
        n11294) );
  nand2_1 U12937 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][26] ), .op(
        n11293) );
  nand2_1 U12938 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][26] ), .op(
        n11292) );
  nand2_1 U12939 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][26] ), .op(
        n11291) );
  and4_1 U12940 ( .ip1(n11294), .ip2(n11293), .ip3(n11292), .ip4(n11291), .op(
        n11321) );
  nand2_1 U12941 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][26] ), .op(
        n11298) );
  nand2_1 U12942 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][26] ), .op(
        n11297) );
  nand2_1 U12943 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][26] ), .op(
        n11296) );
  nand2_1 U12944 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][26] ), .op(
        n11295) );
  and4_1 U12945 ( .ip1(n11298), .ip2(n11297), .ip3(n11296), .ip4(n11295), .op(
        n11320) );
  nand2_1 U12946 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][26] ), .op(
        n11302) );
  nand2_1 U12947 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][26] ), .op(
        n11301) );
  nand2_1 U12948 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][26] ), .op(
        n11300) );
  nand2_1 U12949 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][26] ), .op(
        n11299) );
  nand2_1 U12950 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][26] ), .op(
        n11306) );
  nand2_1 U12951 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][26] ), .op(
        n11305) );
  nand2_1 U12952 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][26] ), .op(
        n11304) );
  nand2_1 U12953 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][26] ), .op(
        n11303) );
  nand2_1 U12954 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][26] ), .op(
        n11310) );
  nand2_1 U12955 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][26] ), .op(
        n11309) );
  nand2_1 U12956 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][26] ), .op(
        n11308) );
  nand2_1 U12957 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][26] ), .op(
        n11307) );
  nand2_1 U12958 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][26] ), .op(
        n11314) );
  nand2_1 U12959 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][26] ), .op(
        n11313) );
  nand2_1 U12960 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][26] ), .op(
        n11312) );
  nand2_1 U12961 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][26] ), .op(
        n11311) );
  mux2_1 U12962 ( .ip1(n19089), .ip2(n11323), .s(n10200), .op(n16333) );
  nand2_1 U12963 ( .ip1(n16333), .ip2(n13520), .op(n11325) );
  nand2_1 U12964 ( .ip1(n13521), .ip2(\pipeline/PC_DX [26]), .op(n11324) );
  nand2_1 U12965 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][26] ), .op(
        n11327) );
  nand2_1 U12966 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][26] ), .op(
        n11326) );
  nand2_1 U12967 ( .ip1(n11327), .ip2(n11326), .op(n11333) );
  nand2_1 U12968 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][26] ), .op(
        n11331) );
  nand2_1 U12969 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][26] ), .op(
        n11330) );
  nand2_1 U12970 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][26] ), .op(
        n11329) );
  nand2_1 U12971 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][26] ), .op(
        n11328) );
  not_ab_or_c_or_d U12972 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][26] ), .ip3(n11333), .ip4(n11332), .op(n11365) );
  nand2_1 U12973 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][26] ), .op(
        n11337) );
  nand2_1 U12974 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][26] ), .op(
        n11336) );
  nand2_1 U12975 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][26] ), .op(
        n11335) );
  nand2_1 U12976 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][26] ), .op(
        n11334) );
  and4_1 U12977 ( .ip1(n11337), .ip2(n11336), .ip3(n11335), .ip4(n11334), .op(
        n11364) );
  nand2_1 U12978 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][26] ), .op(
        n11341) );
  nand2_1 U12979 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][26] ), .op(
        n11340) );
  nand2_1 U12980 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][26] ), .op(
        n11339) );
  nand2_1 U12981 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][26] ), .op(
        n11338) );
  and4_1 U12982 ( .ip1(n11341), .ip2(n11340), .ip3(n11339), .ip4(n11338), .op(
        n11363) );
  nand2_1 U12983 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][26] ), .op(
        n11345) );
  nand2_1 U12984 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][26] ), .op(
        n11344) );
  nand2_1 U12985 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][26] ), .op(
        n11343) );
  nand2_1 U12986 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][26] ), .op(
        n11342) );
  nand2_1 U12987 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][26] ), .op(
        n11349) );
  nand2_1 U12988 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][26] ), .op(
        n11348) );
  nand2_1 U12989 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][26] ), .op(
        n11347) );
  nand2_1 U12990 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][26] ), .op(
        n11346) );
  nand2_1 U12991 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][26] ), .op(
        n11353) );
  nand2_1 U12992 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][26] ), .op(
        n11352) );
  nand2_1 U12993 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][26] ), .op(
        n11351) );
  nand2_1 U12994 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][26] ), .op(
        n11350) );
  nand2_1 U12995 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][26] ), .op(
        n11357) );
  nand2_1 U12996 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][26] ), .op(
        n11356) );
  nand2_1 U12997 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][26] ), .op(
        n11355) );
  nand2_1 U12998 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][26] ), .op(
        n11354) );
  nand2_1 U12999 ( .ip1(n21281), .ip2(n10201), .op(n11370) );
  nor2_1 U13000 ( .ip1(n11367), .ip2(n12836), .op(n11368) );
  nor2_1 U13001 ( .ip1(n12320), .ip2(n11368), .op(n11369) );
  nand2_1 U13002 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [25]), .op(n11373) );
  nand2_1 U13003 ( .ip1(\pipeline/alu_out_WB [25]), .ip2(n17895), .op(n11372)
         );
  nand2_1 U13004 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [25]), .op(
        n11371) );
  nand3_1 U13005 ( .ip1(n11373), .ip2(n11372), .ip3(n11371), .op(n18341) );
  nand2_1 U13006 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][25] ), .op(
        n11375) );
  nand2_1 U13007 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][25] ), .op(
        n11374) );
  nand2_1 U13008 ( .ip1(n11375), .ip2(n11374), .op(n11381) );
  nand2_1 U13009 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][25] ), .op(
        n11379) );
  nand2_1 U13010 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][25] ), .op(
        n11378) );
  nand2_1 U13011 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][25] ), .op(
        n11377) );
  nand2_1 U13012 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][25] ), .op(
        n11376) );
  not_ab_or_c_or_d U13013 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][25] ), .ip3(n11381), .ip4(n11380), .op(n11413) );
  nand2_1 U13014 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][25] ), .op(
        n11385) );
  nand2_1 U13015 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][25] ), .op(
        n11384) );
  nand2_1 U13016 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][25] ), .op(
        n11383) );
  nand2_1 U13017 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][25] ), .op(
        n11382) );
  and4_1 U13018 ( .ip1(n11385), .ip2(n11384), .ip3(n11383), .ip4(n11382), .op(
        n11412) );
  nand2_1 U13019 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][25] ), .op(
        n11389) );
  nand2_1 U13020 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][25] ), .op(
        n11388) );
  nand2_1 U13021 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][25] ), .op(
        n11387) );
  nand2_1 U13022 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][25] ), .op(
        n11386) );
  and4_1 U13023 ( .ip1(n11389), .ip2(n11388), .ip3(n11387), .ip4(n11386), .op(
        n11411) );
  nand2_1 U13024 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][25] ), .op(
        n11393) );
  nand2_1 U13025 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][25] ), .op(
        n11392) );
  nand2_1 U13026 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][25] ), .op(
        n11391) );
  nand2_1 U13027 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][25] ), .op(
        n11390) );
  nand2_1 U13028 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][25] ), .op(
        n11397) );
  nand2_1 U13029 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][25] ), .op(
        n11396) );
  nand2_1 U13030 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][25] ), .op(
        n11395) );
  nand2_1 U13031 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][25] ), .op(
        n11394) );
  nand2_1 U13032 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][25] ), .op(
        n11401) );
  nand2_1 U13033 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][25] ), .op(
        n11400) );
  nand2_1 U13034 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][25] ), .op(
        n11399) );
  nand2_1 U13035 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][25] ), .op(
        n11398) );
  nand2_1 U13036 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][25] ), .op(
        n11405) );
  nand2_1 U13037 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][25] ), .op(
        n11404) );
  nand2_1 U13038 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][25] ), .op(
        n11403) );
  nand2_1 U13039 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][25] ), .op(
        n11402) );
  mux2_1 U13040 ( .ip1(n18341), .ip2(n11414), .s(n10199), .op(n15565) );
  nand2_1 U13041 ( .ip1(n15565), .ip2(n13520), .op(n11416) );
  nand2_1 U13042 ( .ip1(n13521), .ip2(\pipeline/PC_DX [25]), .op(n11415) );
  nand2_1 U13043 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][25] ), .op(
        n11418) );
  nand2_1 U13044 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][25] ), .op(
        n11417) );
  nand2_1 U13045 ( .ip1(n11418), .ip2(n11417), .op(n11424) );
  nand2_1 U13046 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][25] ), .op(
        n11422) );
  nand2_1 U13047 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][25] ), .op(
        n11421) );
  nand2_1 U13048 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][25] ), .op(
        n11420) );
  nand2_1 U13049 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][25] ), .op(
        n11419) );
  not_ab_or_c_or_d U13050 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][25] ), .ip3(n11424), .ip4(n11423), .op(n11456) );
  nand2_1 U13051 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][25] ), .op(
        n11428) );
  nand2_1 U13052 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][25] ), .op(
        n11427) );
  nand2_1 U13053 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][25] ), .op(
        n11426) );
  nand2_1 U13054 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][25] ), .op(
        n11425) );
  and4_1 U13055 ( .ip1(n11428), .ip2(n11427), .ip3(n11426), .ip4(n11425), .op(
        n11455) );
  nand2_1 U13056 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][25] ), .op(
        n11432) );
  nand2_1 U13057 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][25] ), .op(
        n11431) );
  nand2_1 U13058 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][25] ), .op(
        n11430) );
  nand2_1 U13059 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][25] ), .op(
        n11429) );
  and4_1 U13060 ( .ip1(n11432), .ip2(n11431), .ip3(n11430), .ip4(n11429), .op(
        n11454) );
  nand2_1 U13061 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][25] ), .op(
        n11436) );
  nand2_1 U13062 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][25] ), .op(
        n11435) );
  nand2_1 U13063 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][25] ), .op(
        n11434) );
  nand2_1 U13064 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][25] ), .op(
        n11433) );
  nand2_1 U13065 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][25] ), .op(
        n11440) );
  nand2_1 U13066 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][25] ), .op(
        n11439) );
  nand2_1 U13067 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][25] ), .op(
        n11438) );
  nand2_1 U13068 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][25] ), .op(
        n11437) );
  nand2_1 U13069 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][25] ), .op(
        n11444) );
  nand2_1 U13070 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][25] ), .op(
        n11443) );
  nand2_1 U13071 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][25] ), .op(
        n11442) );
  nand2_1 U13072 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][25] ), .op(
        n11441) );
  nand2_1 U13073 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][25] ), .op(
        n11448) );
  nand2_1 U13074 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][25] ), .op(
        n11447) );
  nand2_1 U13075 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][25] ), .op(
        n11446) );
  nand2_1 U13076 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][25] ), .op(
        n11445) );
  nand2_1 U13077 ( .ip1(n21282), .ip2(n10201), .op(n11461) );
  inv_1 U13078 ( .ip(\pipeline/inst_DX [25]), .op(n11458) );
  nor2_1 U13079 ( .ip1(n11458), .ip2(n12836), .op(n11459) );
  nor2_1 U13080 ( .ip1(n12320), .ip2(n11459), .op(n11460) );
  nand2_1 U13081 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [24]), .op(n11464) );
  nand2_1 U13082 ( .ip1(\pipeline/alu_out_WB [24]), .ip2(n17895), .op(n11463)
         );
  nand2_1 U13083 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [24]), .op(
        n11462) );
  nand3_1 U13084 ( .ip1(n11464), .ip2(n11463), .ip3(n11462), .op(n18717) );
  nand2_1 U13085 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][24] ), .op(
        n11466) );
  nand2_1 U13086 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][24] ), .op(
        n11465) );
  nand2_1 U13087 ( .ip1(n11466), .ip2(n11465), .op(n11472) );
  nand2_1 U13088 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][24] ), .op(
        n11470) );
  nand2_1 U13089 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][24] ), .op(
        n11469) );
  nand2_1 U13090 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][24] ), .op(
        n11468) );
  nand2_1 U13091 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][24] ), .op(
        n11467) );
  not_ab_or_c_or_d U13092 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][24] ), .ip3(n11472), .ip4(n11471), .op(n11504) );
  nand2_1 U13093 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][24] ), .op(
        n11476) );
  nand2_1 U13094 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][24] ), .op(
        n11475) );
  nand2_1 U13095 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][24] ), .op(
        n11474) );
  nand2_1 U13096 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][24] ), .op(
        n11473) );
  and4_1 U13097 ( .ip1(n11476), .ip2(n11475), .ip3(n11474), .ip4(n11473), .op(
        n11503) );
  nand2_1 U13098 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][24] ), .op(
        n11480) );
  nand2_1 U13099 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][24] ), .op(
        n11479) );
  nand2_1 U13100 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][24] ), .op(
        n11478) );
  nand2_1 U13101 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][24] ), .op(
        n11477) );
  and4_1 U13102 ( .ip1(n11480), .ip2(n11479), .ip3(n11478), .ip4(n11477), .op(
        n11502) );
  nand2_1 U13103 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][24] ), .op(
        n11484) );
  nand2_1 U13104 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][24] ), .op(
        n11483) );
  nand2_1 U13105 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][24] ), .op(
        n11482) );
  nand2_1 U13106 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][24] ), .op(
        n11481) );
  nand2_1 U13107 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][24] ), .op(
        n11488) );
  nand2_1 U13108 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][24] ), .op(
        n11487) );
  nand2_1 U13109 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][24] ), .op(
        n11486) );
  nand2_1 U13110 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][24] ), .op(
        n11485) );
  nand2_1 U13111 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][24] ), .op(
        n11492) );
  nand2_1 U13112 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][24] ), .op(
        n11491) );
  nand2_1 U13113 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][24] ), .op(
        n11490) );
  nand2_1 U13114 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][24] ), .op(
        n11489) );
  nand2_1 U13115 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][24] ), .op(
        n11496) );
  nand2_1 U13116 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][24] ), .op(
        n11495) );
  nand2_1 U13117 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][24] ), .op(
        n11494) );
  nand2_1 U13118 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][24] ), .op(
        n11493) );
  mux2_1 U13119 ( .ip1(n18717), .ip2(n11505), .s(n10199), .op(n20611) );
  nand2_1 U13120 ( .ip1(n20611), .ip2(n13520), .op(n11507) );
  nand2_1 U13121 ( .ip1(n13521), .ip2(\pipeline/PC_DX [24]), .op(n11506) );
  nand2_1 U13122 ( .ip1(n11507), .ip2(n11506), .op(n11508) );
  nand2_1 U13123 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][24] ), .op(
        n11510) );
  nand2_1 U13124 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][24] ), .op(
        n11509) );
  nand2_1 U13125 ( .ip1(n11510), .ip2(n11509), .op(n11516) );
  nand2_1 U13126 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][24] ), .op(
        n11514) );
  nand2_1 U13127 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][24] ), .op(
        n11513) );
  nand2_1 U13128 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][24] ), .op(
        n11512) );
  nand2_1 U13129 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][24] ), .op(
        n11511) );
  not_ab_or_c_or_d U13130 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][24] ), .ip3(n11516), .ip4(n11515), .op(n11548) );
  nand2_1 U13131 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][24] ), .op(
        n11520) );
  nand2_1 U13132 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][24] ), .op(
        n11519) );
  nand2_1 U13133 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][24] ), .op(
        n11518) );
  nand2_1 U13134 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][24] ), .op(
        n11517) );
  and4_1 U13135 ( .ip1(n11520), .ip2(n11519), .ip3(n11518), .ip4(n11517), .op(
        n11547) );
  nand2_1 U13136 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][24] ), .op(
        n11524) );
  nand2_1 U13137 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][24] ), .op(
        n11523) );
  nand2_1 U13138 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][24] ), .op(
        n11522) );
  nand2_1 U13139 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][24] ), .op(
        n11521) );
  and4_1 U13140 ( .ip1(n11524), .ip2(n11523), .ip3(n11522), .ip4(n11521), .op(
        n11546) );
  nand2_1 U13141 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][24] ), .op(
        n11528) );
  nand2_1 U13142 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][24] ), .op(
        n11527) );
  nand2_1 U13143 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][24] ), .op(
        n11526) );
  nand2_1 U13144 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][24] ), .op(
        n11525) );
  nand2_1 U13145 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][24] ), .op(
        n11532) );
  nand2_1 U13146 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][24] ), .op(
        n11531) );
  nand2_1 U13147 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][24] ), .op(
        n11530) );
  nand2_1 U13148 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][24] ), .op(
        n11529) );
  nand2_1 U13149 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][24] ), .op(
        n11536) );
  nand2_1 U13150 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][24] ), .op(
        n11535) );
  nand2_1 U13151 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][24] ), .op(
        n11534) );
  nand2_1 U13152 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][24] ), .op(
        n11533) );
  nand2_1 U13153 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][24] ), .op(
        n11540) );
  nand2_1 U13154 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][24] ), .op(
        n11539) );
  nand2_1 U13155 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][24] ), .op(
        n11538) );
  nand2_1 U13156 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][24] ), .op(
        n11537) );
  buf_4 U13157 ( .ip(n13063), .op(n13315) );
  buf_4 U13158 ( .ip(n13315), .op(n12683) );
  mux2_1 U13159 ( .ip1(n18717), .ip2(n11549), .s(n12683), .op(n21278) );
  nand2_1 U13160 ( .ip1(n21278), .ip2(n10201), .op(n11552) );
  nor2_1 U13161 ( .ip1(n12837), .ip2(n12836), .op(n11550) );
  nor2_1 U13162 ( .ip1(n12320), .ip2(n11550), .op(n11551) );
  nand2_1 U13163 ( .ip1(n11552), .ip2(n11551), .op(n18731) );
  nor2_1 U13164 ( .ip1(n13656), .ip2(n18731), .op(n11553) );
  nor2_1 U13165 ( .ip1(n11938), .ip2(n11553), .op(n11554) );
  nand2_1 U13166 ( .ip1(n11943), .ip2(n11554), .op(n11926) );
  nand2_1 U13167 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [30]), .op(n11557) );
  nand2_1 U13168 ( .ip1(\pipeline/alu_out_WB [30]), .ip2(n17895), .op(n11556)
         );
  nand2_1 U13169 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [30]), .op(
        n11555) );
  nand3_1 U13170 ( .ip1(n11557), .ip2(n11556), .ip3(n11555), .op(n18867) );
  nand2_1 U13171 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][30] ), .op(
        n11559) );
  nand2_1 U13172 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][30] ), .op(
        n11558) );
  nand2_1 U13173 ( .ip1(n11559), .ip2(n11558), .op(n11565) );
  nand2_1 U13174 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][30] ), .op(
        n11563) );
  nand2_1 U13175 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][30] ), .op(
        n11562) );
  nand2_1 U13176 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][30] ), .op(
        n11561) );
  nand2_1 U13177 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][30] ), .op(
        n11560) );
  not_ab_or_c_or_d U13178 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][30] ), .ip3(n11565), .ip4(n11564), .op(n11597) );
  nand2_1 U13179 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][30] ), .op(
        n11569) );
  nand2_1 U13180 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][30] ), .op(
        n11568) );
  nand2_1 U13181 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][30] ), .op(
        n11567) );
  nand2_1 U13182 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][30] ), .op(
        n11566) );
  and4_1 U13183 ( .ip1(n11569), .ip2(n11568), .ip3(n11567), .ip4(n11566), .op(
        n11596) );
  nand2_1 U13184 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][30] ), .op(
        n11573) );
  nand2_1 U13185 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][30] ), .op(
        n11572) );
  nand2_1 U13186 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][30] ), .op(
        n11571) );
  nand2_1 U13187 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][30] ), .op(
        n11570) );
  and4_1 U13188 ( .ip1(n11573), .ip2(n11572), .ip3(n11571), .ip4(n11570), .op(
        n11595) );
  nand2_1 U13189 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][30] ), .op(
        n11577) );
  nand2_1 U13190 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][30] ), .op(
        n11576) );
  nand2_1 U13191 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][30] ), .op(
        n11575) );
  nand2_1 U13192 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][30] ), .op(
        n11574) );
  nand2_1 U13193 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][30] ), .op(
        n11581) );
  nand2_1 U13194 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][30] ), .op(
        n11580) );
  nand2_1 U13195 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][30] ), .op(
        n11579) );
  nand2_1 U13196 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][30] ), .op(
        n11578) );
  nand2_1 U13197 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][30] ), .op(
        n11585) );
  nand2_1 U13198 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][30] ), .op(
        n11584) );
  nand2_1 U13199 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][30] ), .op(
        n11583) );
  nand2_1 U13200 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][30] ), .op(
        n11582) );
  nand2_1 U13201 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][30] ), .op(
        n11589) );
  nand2_1 U13202 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][30] ), .op(
        n11588) );
  nand2_1 U13203 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][30] ), .op(
        n11587) );
  nand2_1 U13204 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][30] ), .op(
        n11586) );
  mux2_1 U13205 ( .ip1(n18867), .ip2(n11598), .s(n10199), .op(n21645) );
  nand2_1 U13206 ( .ip1(n21645), .ip2(n13520), .op(n11600) );
  nand2_1 U13207 ( .ip1(n13521), .ip2(\pipeline/PC_DX [30]), .op(n11599) );
  nand2_1 U13208 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][30] ), .op(
        n11602) );
  nand2_1 U13209 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][30] ), .op(
        n11601) );
  nand2_1 U13210 ( .ip1(n11602), .ip2(n11601), .op(n11608) );
  nand2_1 U13211 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][30] ), .op(
        n11606) );
  nand2_1 U13212 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][30] ), .op(
        n11605) );
  nand2_1 U13213 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][30] ), .op(
        n11604) );
  nand2_1 U13214 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][30] ), .op(
        n11603) );
  not_ab_or_c_or_d U13215 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][30] ), .ip3(n11608), .ip4(n11607), .op(n11640) );
  nand2_1 U13216 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][30] ), .op(
        n11612) );
  nand2_1 U13217 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][30] ), .op(
        n11611) );
  nand2_1 U13218 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][30] ), .op(
        n11610) );
  nand2_1 U13219 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][30] ), .op(
        n11609) );
  and4_1 U13220 ( .ip1(n11612), .ip2(n11611), .ip3(n11610), .ip4(n11609), .op(
        n11639) );
  nand2_1 U13221 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][30] ), .op(
        n11616) );
  nand2_1 U13222 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][30] ), .op(
        n11615) );
  nand2_1 U13223 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][30] ), .op(
        n11614) );
  nand2_1 U13224 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][30] ), .op(
        n11613) );
  and4_1 U13225 ( .ip1(n11616), .ip2(n11615), .ip3(n11614), .ip4(n11613), .op(
        n11638) );
  nand2_1 U13226 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][30] ), .op(
        n11620) );
  nand2_1 U13227 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][30] ), .op(
        n11619) );
  nand2_1 U13228 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][30] ), .op(
        n11618) );
  nand2_1 U13229 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][30] ), .op(
        n11617) );
  nand2_1 U13230 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][30] ), .op(
        n11624) );
  nand2_1 U13231 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][30] ), .op(
        n11623) );
  nand2_1 U13232 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][30] ), .op(
        n11622) );
  nand2_1 U13233 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][30] ), .op(
        n11621) );
  nand2_1 U13234 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][30] ), .op(
        n11628) );
  nand2_1 U13235 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][30] ), .op(
        n11627) );
  nand2_1 U13236 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][30] ), .op(
        n11626) );
  nand2_1 U13237 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][30] ), .op(
        n11625) );
  nand2_1 U13238 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][30] ), .op(
        n11632) );
  nand2_1 U13239 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][30] ), .op(
        n11631) );
  nand2_1 U13240 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][30] ), .op(
        n11630) );
  nand2_1 U13241 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][30] ), .op(
        n11629) );
  inv_1 U13242 ( .ip(\pipeline/inst_DX [30]), .op(n15308) );
  nor2_1 U13243 ( .ip1(n15308), .ip2(n12836), .op(n11642) );
  nor2_1 U13244 ( .ip1(n12320), .ip2(n11642), .op(n11643) );
  nor2_1 U13245 ( .ip1(n10181), .ip2(n17102), .op(n11737) );
  nand2_1 U13246 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [31]), .op(n11647) );
  nand2_1 U13247 ( .ip1(\pipeline/alu_out_WB [31]), .ip2(n17895), .op(n11646)
         );
  nand2_1 U13248 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [31]), .op(
        n11645) );
  nand3_1 U13249 ( .ip1(n11647), .ip2(n11646), .ip3(n11645), .op(n21584) );
  nand2_1 U13250 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][31] ), .op(
        n11649) );
  nand2_1 U13251 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][31] ), .op(
        n11648) );
  nand2_1 U13252 ( .ip1(n11649), .ip2(n11648), .op(n11655) );
  nand2_1 U13253 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][31] ), .op(
        n11653) );
  nand2_1 U13254 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][31] ), .op(
        n11652) );
  nand2_1 U13255 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][31] ), .op(
        n11651) );
  nand2_1 U13256 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][31] ), .op(
        n11650) );
  not_ab_or_c_or_d U13257 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][31] ), .ip3(n11655), .ip4(n11654), .op(n11687) );
  nand2_1 U13258 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][31] ), .op(
        n11659) );
  nand2_1 U13259 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][31] ), .op(
        n11658) );
  nand2_1 U13260 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][31] ), .op(
        n11657) );
  nand2_1 U13261 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][31] ), .op(
        n11656) );
  and4_1 U13262 ( .ip1(n11659), .ip2(n11658), .ip3(n11657), .ip4(n11656), .op(
        n11686) );
  nand2_1 U13263 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][31] ), .op(
        n11663) );
  nand2_1 U13264 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][31] ), .op(
        n11662) );
  nand2_1 U13265 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][31] ), .op(
        n11661) );
  nand2_1 U13266 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][31] ), .op(
        n11660) );
  and4_1 U13267 ( .ip1(n11663), .ip2(n11662), .ip3(n11661), .ip4(n11660), .op(
        n11685) );
  nand2_1 U13268 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][31] ), .op(
        n11667) );
  nand2_1 U13269 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][31] ), .op(
        n11666) );
  nand2_1 U13270 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][31] ), .op(
        n11665) );
  nand2_1 U13271 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][31] ), .op(
        n11664) );
  nand2_1 U13272 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][31] ), .op(
        n11671) );
  nand2_1 U13273 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][31] ), .op(
        n11670) );
  nand2_1 U13274 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][31] ), .op(
        n11669) );
  nand2_1 U13275 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][31] ), .op(
        n11668) );
  nand2_1 U13276 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][31] ), .op(
        n11675) );
  nand2_1 U13277 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][31] ), .op(
        n11674) );
  nand2_1 U13278 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][31] ), .op(
        n11673) );
  nand2_1 U13279 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][31] ), .op(
        n11672) );
  nand2_1 U13280 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][31] ), .op(
        n11679) );
  nand2_1 U13281 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][31] ), .op(
        n11678) );
  nand2_1 U13282 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][31] ), .op(
        n11677) );
  nand2_1 U13283 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][31] ), .op(
        n11676) );
  mux2_1 U13284 ( .ip1(n21584), .ip2(n11688), .s(n10199), .op(n14594) );
  nand2_1 U13285 ( .ip1(n14594), .ip2(n13520), .op(n11690) );
  nand2_1 U13286 ( .ip1(n13521), .ip2(\pipeline/PC_DX [31]), .op(n11689) );
  nand2_1 U13287 ( .ip1(n11690), .ip2(n11689), .op(n11934) );
  nand2_1 U13288 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][31] ), .op(
        n11693) );
  nand2_1 U13289 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][31] ), .op(
        n11692) );
  nand2_1 U13290 ( .ip1(n11693), .ip2(n11692), .op(n11699) );
  nand2_1 U13291 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][31] ), .op(
        n11697) );
  nand2_1 U13292 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][31] ), .op(
        n11696) );
  nand2_1 U13293 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][31] ), .op(
        n11695) );
  nand2_1 U13294 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][31] ), .op(
        n11694) );
  not_ab_or_c_or_d U13295 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][31] ), .ip3(n11699), .ip4(n11698), .op(n11731) );
  nand2_1 U13296 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][31] ), .op(
        n11703) );
  nand2_1 U13297 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][31] ), .op(
        n11702) );
  nand2_1 U13298 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][31] ), .op(
        n11701) );
  nand2_1 U13299 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][31] ), .op(
        n11700) );
  and4_1 U13300 ( .ip1(n11703), .ip2(n11702), .ip3(n11701), .ip4(n11700), .op(
        n11730) );
  nand2_1 U13301 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][31] ), .op(
        n11707) );
  nand2_1 U13302 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][31] ), .op(
        n11706) );
  nand2_1 U13303 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][31] ), .op(
        n11705) );
  nand2_1 U13304 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][31] ), .op(
        n11704) );
  and4_1 U13305 ( .ip1(n11707), .ip2(n11706), .ip3(n11705), .ip4(n11704), .op(
        n11729) );
  nand2_1 U13306 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][31] ), .op(
        n11711) );
  nand2_1 U13307 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][31] ), .op(
        n11710) );
  nand2_1 U13308 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][31] ), .op(
        n11709) );
  nand2_1 U13309 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][31] ), .op(
        n11708) );
  nand2_1 U13310 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][31] ), .op(
        n11715) );
  nand2_1 U13311 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][31] ), .op(
        n11714) );
  nand2_1 U13312 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][31] ), .op(
        n11713) );
  nand2_1 U13313 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][31] ), .op(
        n11712) );
  nand2_1 U13314 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][31] ), .op(
        n11719) );
  nand2_1 U13315 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][31] ), .op(
        n11718) );
  nand2_1 U13316 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][31] ), .op(
        n11717) );
  nand2_1 U13317 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][31] ), .op(
        n11716) );
  nand2_1 U13318 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][31] ), .op(
        n11723) );
  nand2_1 U13319 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][31] ), .op(
        n11722) );
  nand2_1 U13320 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][31] ), .op(
        n11721) );
  nand2_1 U13321 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][31] ), .op(
        n11720) );
  nand2_1 U13322 ( .ip1(n11732), .ip2(n13315), .op(n11733) );
  inv_1 U13323 ( .ip(n13209), .op(n13220) );
  nand2_1 U13324 ( .ip1(\pipeline/imm[31] ), .ip2(n13220), .op(n11735) );
  nand2_2 U13325 ( .ip1(n11736), .ip2(n11735), .op(n20903) );
  nor2_1 U13326 ( .ip1(n11737), .ip2(n13978), .op(n11932) );
  nand2_1 U13327 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [29]), .op(n11740) );
  nand2_1 U13328 ( .ip1(\pipeline/alu_out_WB [29]), .ip2(n17895), .op(n11739)
         );
  nand2_1 U13329 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [29]), .op(
        n11738) );
  nand3_1 U13330 ( .ip1(n11740), .ip2(n11739), .ip3(n11738), .op(n18040) );
  nand2_1 U13331 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][29] ), .op(
        n11742) );
  nand2_1 U13332 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][29] ), .op(
        n11741) );
  nand2_1 U13333 ( .ip1(n11742), .ip2(n11741), .op(n11748) );
  nand2_1 U13334 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][29] ), .op(
        n11746) );
  nand2_1 U13335 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][29] ), .op(
        n11745) );
  nand2_1 U13336 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][29] ), .op(
        n11744) );
  nand2_1 U13337 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][29] ), .op(
        n11743) );
  not_ab_or_c_or_d U13338 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][29] ), .ip3(n11748), .ip4(n11747), .op(n11780) );
  nand2_1 U13339 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][29] ), .op(
        n11752) );
  nand2_1 U13340 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][29] ), .op(
        n11751) );
  nand2_1 U13341 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][29] ), .op(
        n11750) );
  nand2_1 U13342 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][29] ), .op(
        n11749) );
  and4_1 U13343 ( .ip1(n11752), .ip2(n11751), .ip3(n11750), .ip4(n11749), .op(
        n11779) );
  nand2_1 U13344 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][29] ), .op(
        n11756) );
  nand2_1 U13345 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][29] ), .op(
        n11755) );
  nand2_1 U13346 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][29] ), .op(
        n11754) );
  nand2_1 U13347 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][29] ), .op(
        n11753) );
  and4_1 U13348 ( .ip1(n11756), .ip2(n11755), .ip3(n11754), .ip4(n11753), .op(
        n11778) );
  nand2_1 U13349 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][29] ), .op(
        n11760) );
  nand2_1 U13350 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][29] ), .op(
        n11759) );
  nand2_1 U13351 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][29] ), .op(
        n11758) );
  nand2_1 U13352 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][29] ), .op(
        n11757) );
  nand2_1 U13353 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][29] ), .op(
        n11764) );
  nand2_1 U13354 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][29] ), .op(
        n11763) );
  nand2_1 U13355 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][29] ), .op(
        n11762) );
  nand2_1 U13356 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][29] ), .op(
        n11761) );
  nand2_1 U13357 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][29] ), .op(
        n11768) );
  nand2_1 U13358 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][29] ), .op(
        n11767) );
  nand2_1 U13359 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][29] ), .op(
        n11766) );
  nand2_1 U13360 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][29] ), .op(
        n11765) );
  nand2_1 U13361 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][29] ), .op(
        n11772) );
  nand2_1 U13362 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][29] ), .op(
        n11771) );
  nand2_1 U13363 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][29] ), .op(
        n11770) );
  nand2_1 U13364 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][29] ), .op(
        n11769) );
  mux2_1 U13365 ( .ip1(n18040), .ip2(n11781), .s(n10199), .op(n20650) );
  nand2_1 U13366 ( .ip1(n20650), .ip2(n13520), .op(n11783) );
  nand2_1 U13367 ( .ip1(\pipeline/PC_DX [29]), .ip2(n13521), .op(n11782) );
  nand2_1 U13368 ( .ip1(n11783), .ip2(n11782), .op(n13599) );
  nand2_1 U13369 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][29] ), .op(
        n11786) );
  nand2_1 U13370 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][29] ), .op(
        n11785) );
  nand2_1 U13371 ( .ip1(n11786), .ip2(n11785), .op(n11792) );
  nand2_1 U13372 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][29] ), .op(
        n11790) );
  nand2_1 U13373 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][29] ), .op(
        n11789) );
  nand2_1 U13374 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][29] ), .op(
        n11788) );
  nand2_1 U13375 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][29] ), .op(
        n11787) );
  not_ab_or_c_or_d U13376 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][29] ), .ip3(n11792), .ip4(n11791), .op(n11824) );
  nand2_1 U13377 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][29] ), .op(
        n11796) );
  nand2_1 U13378 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][29] ), .op(
        n11795) );
  nand2_1 U13379 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][29] ), .op(
        n11794) );
  nand2_1 U13380 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][29] ), .op(
        n11793) );
  and4_1 U13381 ( .ip1(n11796), .ip2(n11795), .ip3(n11794), .ip4(n11793), .op(
        n11823) );
  nand2_1 U13382 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][29] ), .op(
        n11800) );
  nand2_1 U13383 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][29] ), .op(
        n11799) );
  nand2_1 U13384 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][29] ), .op(
        n11798) );
  nand2_1 U13385 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][29] ), .op(
        n11797) );
  and4_1 U13386 ( .ip1(n11800), .ip2(n11799), .ip3(n11798), .ip4(n11797), .op(
        n11822) );
  nand2_1 U13387 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][29] ), .op(
        n11804) );
  nand2_1 U13388 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][29] ), .op(
        n11803) );
  nand2_1 U13389 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][29] ), .op(
        n11802) );
  nand2_1 U13390 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][29] ), .op(
        n11801) );
  nand2_1 U13391 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][29] ), .op(
        n11808) );
  nand2_1 U13392 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][29] ), .op(
        n11807) );
  nand2_1 U13393 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][29] ), .op(
        n11806) );
  nand2_1 U13394 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][29] ), .op(
        n11805) );
  nand2_1 U13395 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][29] ), .op(
        n11812) );
  nand2_1 U13396 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][29] ), .op(
        n11811) );
  nand2_1 U13397 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][29] ), .op(
        n11810) );
  nand2_1 U13398 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][29] ), .op(
        n11809) );
  nand2_1 U13399 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][29] ), .op(
        n11816) );
  nand2_1 U13400 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][29] ), .op(
        n11815) );
  nand2_1 U13401 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][29] ), .op(
        n11814) );
  nand2_1 U13402 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][29] ), .op(
        n11813) );
  inv_1 U13403 ( .ip(\pipeline/inst_DX [29]), .op(n22121) );
  nor2_1 U13404 ( .ip1(n22121), .ip2(n12836), .op(n11828) );
  nor2_1 U13405 ( .ip1(n12320), .ip2(n11828), .op(n11829) );
  nand2_1 U13406 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [28]), .op(n11833) );
  nand2_1 U13407 ( .ip1(\pipeline/alu_out_WB [28]), .ip2(n17895), .op(n11832)
         );
  nand2_1 U13408 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [28]), .op(
        n11831) );
  nand3_1 U13409 ( .ip1(n11833), .ip2(n11832), .ip3(n11831), .op(n19032) );
  nand2_1 U13410 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][28] ), .op(
        n11835) );
  nand2_1 U13411 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][28] ), .op(
        n11834) );
  nand2_1 U13412 ( .ip1(n11835), .ip2(n11834), .op(n11841) );
  nand2_1 U13413 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][28] ), .op(
        n11839) );
  nand2_1 U13414 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][28] ), .op(
        n11838) );
  nand2_1 U13415 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][28] ), .op(
        n11837) );
  nand2_1 U13416 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][28] ), .op(
        n11836) );
  not_ab_or_c_or_d U13417 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][28] ), .ip3(n11841), .ip4(n11840), .op(n11873) );
  nand2_1 U13418 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][28] ), .op(
        n11845) );
  nand2_1 U13419 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][28] ), .op(
        n11844) );
  nand2_1 U13420 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][28] ), .op(
        n11843) );
  nand2_1 U13421 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][28] ), .op(
        n11842) );
  and4_1 U13422 ( .ip1(n11845), .ip2(n11844), .ip3(n11843), .ip4(n11842), .op(
        n11872) );
  nand2_1 U13423 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][28] ), .op(
        n11849) );
  nand2_1 U13424 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][28] ), .op(
        n11848) );
  nand2_1 U13425 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][28] ), .op(
        n11847) );
  nand2_1 U13426 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][28] ), .op(
        n11846) );
  and4_1 U13427 ( .ip1(n11849), .ip2(n11848), .ip3(n11847), .ip4(n11846), .op(
        n11871) );
  nand2_1 U13428 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][28] ), .op(
        n11853) );
  nand2_1 U13429 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][28] ), .op(
        n11852) );
  nand2_1 U13430 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][28] ), .op(
        n11851) );
  nand2_1 U13431 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][28] ), .op(
        n11850) );
  nand2_1 U13432 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][28] ), .op(
        n11857) );
  nand2_1 U13433 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][28] ), .op(
        n11856) );
  nand2_1 U13434 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][28] ), .op(
        n11855) );
  nand2_1 U13435 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][28] ), .op(
        n11854) );
  nand2_1 U13436 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][28] ), .op(
        n11861) );
  nand2_1 U13437 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][28] ), .op(
        n11860) );
  nand2_1 U13438 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][28] ), .op(
        n11859) );
  nand2_1 U13439 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][28] ), .op(
        n11858) );
  nand2_1 U13440 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][28] ), .op(
        n11865) );
  nand2_1 U13441 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][28] ), .op(
        n11864) );
  nand2_1 U13442 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][28] ), .op(
        n11863) );
  nand2_1 U13443 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][28] ), .op(
        n11862) );
  mux2_1 U13444 ( .ip1(n19032), .ip2(n11874), .s(n10200), .op(n20646) );
  nand2_1 U13445 ( .ip1(n20646), .ip2(n13520), .op(n11876) );
  nand2_1 U13446 ( .ip1(n13521), .ip2(\pipeline/PC_DX [28]), .op(n11875) );
  nand2_1 U13447 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][28] ), .op(
        n11879) );
  nand2_1 U13448 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][28] ), .op(
        n11878) );
  nand2_1 U13449 ( .ip1(n11879), .ip2(n11878), .op(n11885) );
  nand2_1 U13450 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][28] ), .op(
        n11883) );
  nand2_1 U13451 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][28] ), .op(
        n11882) );
  nand2_1 U13452 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][28] ), .op(
        n11881) );
  nand2_1 U13453 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][28] ), .op(
        n11880) );
  not_ab_or_c_or_d U13454 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][28] ), .ip3(n11885), .ip4(n11884), .op(n11917) );
  nand2_1 U13455 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][28] ), .op(
        n11889) );
  nand2_1 U13456 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][28] ), .op(
        n11888) );
  nand2_1 U13457 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][28] ), .op(
        n11887) );
  nand2_1 U13458 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][28] ), .op(
        n11886) );
  and4_1 U13459 ( .ip1(n11889), .ip2(n11888), .ip3(n11887), .ip4(n11886), .op(
        n11916) );
  nand2_1 U13460 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][28] ), .op(
        n11893) );
  nand2_1 U13461 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][28] ), .op(
        n11892) );
  nand2_1 U13462 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][28] ), .op(
        n11891) );
  nand2_1 U13463 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][28] ), .op(
        n11890) );
  and4_1 U13464 ( .ip1(n11893), .ip2(n11892), .ip3(n11891), .ip4(n11890), .op(
        n11915) );
  nand2_1 U13465 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][28] ), .op(
        n11897) );
  nand2_1 U13466 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][28] ), .op(
        n11896) );
  nand2_1 U13467 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][28] ), .op(
        n11895) );
  nand2_1 U13468 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][28] ), .op(
        n11894) );
  nand2_1 U13469 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][28] ), .op(
        n11901) );
  nand2_1 U13470 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][28] ), .op(
        n11900) );
  nand2_1 U13471 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][28] ), .op(
        n11899) );
  nand2_1 U13472 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][28] ), .op(
        n11898) );
  nand2_1 U13473 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][28] ), .op(
        n11905) );
  nand2_1 U13474 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][28] ), .op(
        n11904) );
  nand2_1 U13475 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][28] ), .op(
        n11903) );
  nand2_1 U13476 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][28] ), .op(
        n11902) );
  nand2_1 U13477 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][28] ), .op(
        n11909) );
  nand2_1 U13478 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][28] ), .op(
        n11908) );
  nand2_1 U13479 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][28] ), .op(
        n11907) );
  nand2_1 U13480 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][28] ), .op(
        n11906) );
  nor2_1 U13481 ( .ip1(n22120), .ip2(n12836), .op(n11921) );
  nor2_1 U13482 ( .ip1(n12320), .ip2(n11921), .op(n11922) );
  nor2_1 U13483 ( .ip1(n10180), .ip2(n19069), .op(n11924) );
  nor2_1 U13484 ( .ip1(n11928), .ip2(n11924), .op(n11925) );
  nand2_1 U13485 ( .ip1(n11932), .ip2(n11925), .op(n11950) );
  nor2_1 U13486 ( .ip1(n11926), .ip2(n11950), .op(n13570) );
  nand2_1 U13487 ( .ip1(n10180), .ip2(n19069), .op(n11929) );
  or2_1 U13488 ( .ip1(n11929), .ip2(n11928), .op(n11931) );
  nand2_1 U13489 ( .ip1(n10191), .ip2(n18920), .op(n11930) );
  inv_1 U13490 ( .ip(n11934), .op(n13596) );
  nand2_1 U13491 ( .ip1(n13596), .ip2(n20903), .op(n13995) );
  nand2_1 U13492 ( .ip1(n10181), .ip2(n17102), .op(n11935) );
  or2_1 U13493 ( .ip1(n11935), .ip2(n13978), .op(n11936) );
  nand2_1 U13494 ( .ip1(n16533), .ip2(n13601), .op(n11948) );
  nand2_1 U13495 ( .ip1(n10178), .ip2(n16935), .op(n11946) );
  or2_1 U13496 ( .ip1(n11946), .ip2(n11945), .op(n11947) );
  nand2_1 U13497 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [15]), .op(n11958) );
  nand2_1 U13498 ( .ip1(\pipeline/alu_out_WB [15]), .ip2(n17895), .op(n11957)
         );
  nand2_1 U13499 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [15]), .op(
        n11956) );
  nand3_1 U13500 ( .ip1(n11958), .ip2(n11957), .ip3(n11956), .op(n18283) );
  nand2_1 U13501 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][15] ), .op(
        n11960) );
  nand2_1 U13502 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][15] ), .op(
        n11959) );
  nand2_1 U13503 ( .ip1(n11960), .ip2(n11959), .op(n11966) );
  nand2_1 U13504 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][15] ), .op(
        n11964) );
  nand2_1 U13505 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][15] ), .op(
        n11963) );
  nand2_1 U13506 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][15] ), .op(
        n11962) );
  nand2_1 U13507 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][15] ), .op(
        n11961) );
  not_ab_or_c_or_d U13508 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][15] ), .ip3(n11966), .ip4(n11965), .op(n11998) );
  nand2_1 U13509 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][15] ), .op(
        n11970) );
  nand2_1 U13510 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][15] ), .op(
        n11969) );
  nand2_1 U13511 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][15] ), .op(
        n11968) );
  nand2_1 U13512 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][15] ), .op(
        n11967) );
  and4_1 U13513 ( .ip1(n11970), .ip2(n11969), .ip3(n11968), .ip4(n11967), .op(
        n11997) );
  nand2_1 U13514 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][15] ), .op(
        n11974) );
  nand2_1 U13515 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][15] ), .op(
        n11973) );
  nand2_1 U13516 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][15] ), .op(
        n11972) );
  nand2_1 U13517 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][15] ), .op(
        n11971) );
  and4_1 U13518 ( .ip1(n11974), .ip2(n11973), .ip3(n11972), .ip4(n11971), .op(
        n11996) );
  nand2_1 U13519 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][15] ), .op(
        n11978) );
  nand2_1 U13520 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][15] ), .op(
        n11977) );
  nand2_1 U13521 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][15] ), .op(
        n11976) );
  nand2_1 U13522 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][15] ), .op(
        n11975) );
  nand2_1 U13523 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][15] ), .op(
        n11982) );
  nand2_1 U13524 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][15] ), .op(
        n11981) );
  nand2_1 U13525 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][15] ), .op(
        n11980) );
  nand2_1 U13526 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][15] ), .op(
        n11979) );
  nand2_1 U13527 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][15] ), .op(
        n11986) );
  nand2_1 U13528 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][15] ), .op(
        n11985) );
  nand2_1 U13529 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][15] ), .op(
        n11984) );
  nand2_1 U13530 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][15] ), .op(
        n11983) );
  nand2_1 U13531 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][15] ), .op(
        n11990) );
  nand2_1 U13532 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][15] ), .op(
        n11989) );
  nand2_1 U13533 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][15] ), .op(
        n11988) );
  nand2_1 U13534 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][15] ), .op(
        n11987) );
  mux2_1 U13535 ( .ip1(n18283), .ip2(n12000), .s(n10200), .op(n20426) );
  nand2_1 U13536 ( .ip1(n20426), .ip2(n13520), .op(n12002) );
  nand2_1 U13537 ( .ip1(n13521), .ip2(\pipeline/PC_DX [15]), .op(n12001) );
  nand2_1 U13538 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][15] ), .op(
        n12004) );
  nand2_1 U13539 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][15] ), .op(
        n12003) );
  nand2_1 U13540 ( .ip1(n12004), .ip2(n12003), .op(n12010) );
  nand2_1 U13541 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][15] ), .op(
        n12008) );
  nand2_1 U13542 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][15] ), .op(
        n12007) );
  nand2_1 U13543 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][15] ), .op(
        n12006) );
  nand2_1 U13544 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][15] ), .op(
        n12005) );
  not_ab_or_c_or_d U13545 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][15] ), .ip3(n12010), .ip4(n12009), .op(n12042) );
  nand2_1 U13546 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][15] ), .op(
        n12014) );
  nand2_1 U13547 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][15] ), .op(
        n12013) );
  nand2_1 U13548 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][15] ), .op(
        n12012) );
  nand2_1 U13549 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][15] ), .op(
        n12011) );
  and4_1 U13550 ( .ip1(n12014), .ip2(n12013), .ip3(n12012), .ip4(n12011), .op(
        n12041) );
  nand2_1 U13551 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][15] ), .op(
        n12018) );
  nand2_1 U13552 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][15] ), .op(
        n12017) );
  nand2_1 U13553 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][15] ), .op(
        n12016) );
  nand2_1 U13554 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][15] ), .op(
        n12015) );
  and4_1 U13555 ( .ip1(n12018), .ip2(n12017), .ip3(n12016), .ip4(n12015), .op(
        n12040) );
  nand2_1 U13556 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][15] ), .op(
        n12022) );
  nand2_1 U13557 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][15] ), .op(
        n12021) );
  nand2_1 U13558 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][15] ), .op(
        n12020) );
  nand2_1 U13559 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][15] ), .op(
        n12019) );
  nand2_1 U13560 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][15] ), .op(
        n12026) );
  nand2_1 U13561 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][15] ), .op(
        n12025) );
  nand2_1 U13562 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][15] ), .op(
        n12024) );
  nand2_1 U13563 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][15] ), .op(
        n12023) );
  nand2_1 U13564 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][15] ), .op(
        n12030) );
  nand2_1 U13565 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][15] ), .op(
        n12029) );
  nand2_1 U13566 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][15] ), .op(
        n12028) );
  nand2_1 U13567 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][15] ), .op(
        n12027) );
  nand2_1 U13568 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][15] ), .op(
        n12034) );
  nand2_1 U13569 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][15] ), .op(
        n12033) );
  nand2_1 U13570 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][15] ), .op(
        n12032) );
  nand2_1 U13571 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][15] ), .op(
        n12031) );
  nor2_1 U13572 ( .ip1(n16028), .ip2(n12836), .op(n12044) );
  nor2_1 U13573 ( .ip1(n12320), .ip2(n12044), .op(n12045) );
  nand2_1 U13574 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [14]), .op(n12049) );
  nand2_1 U13575 ( .ip1(\pipeline/alu_out_WB [14]), .ip2(n17895), .op(n12048)
         );
  nand2_1 U13576 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [14]), .op(
        n12047) );
  nand3_1 U13577 ( .ip1(n12049), .ip2(n12048), .ip3(n12047), .op(n19330) );
  nand2_1 U13578 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][14] ), .op(
        n12051) );
  nand2_1 U13579 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][14] ), .op(
        n12050) );
  nand2_1 U13580 ( .ip1(n12051), .ip2(n12050), .op(n12057) );
  nand2_1 U13581 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][14] ), .op(
        n12055) );
  nand2_1 U13582 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][14] ), .op(
        n12054) );
  nand2_1 U13583 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][14] ), .op(
        n12053) );
  nand2_1 U13584 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][14] ), .op(
        n12052) );
  not_ab_or_c_or_d U13585 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][14] ), .ip3(n12057), .ip4(n12056), .op(n12089) );
  nand2_1 U13586 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][14] ), .op(
        n12061) );
  nand2_1 U13587 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][14] ), .op(
        n12060) );
  nand2_1 U13588 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][14] ), .op(
        n12059) );
  nand2_1 U13589 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][14] ), .op(
        n12058) );
  and4_1 U13590 ( .ip1(n12061), .ip2(n12060), .ip3(n12059), .ip4(n12058), .op(
        n12088) );
  nand2_1 U13591 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][14] ), .op(
        n12065) );
  nand2_1 U13592 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][14] ), .op(
        n12064) );
  nand2_1 U13593 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][14] ), .op(
        n12063) );
  nand2_1 U13594 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][14] ), .op(
        n12062) );
  and4_1 U13595 ( .ip1(n12065), .ip2(n12064), .ip3(n12063), .ip4(n12062), .op(
        n12087) );
  nand2_1 U13596 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][14] ), .op(
        n12069) );
  nand2_1 U13597 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][14] ), .op(
        n12068) );
  nand2_1 U13598 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][14] ), .op(
        n12067) );
  nand2_1 U13599 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][14] ), .op(
        n12066) );
  nand2_1 U13600 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][14] ), .op(
        n12073) );
  nand2_1 U13601 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][14] ), .op(
        n12072) );
  nand2_1 U13602 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][14] ), .op(
        n12071) );
  nand2_1 U13603 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][14] ), .op(
        n12070) );
  nand2_1 U13604 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][14] ), .op(
        n12077) );
  nand2_1 U13605 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][14] ), .op(
        n12076) );
  nand2_1 U13606 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][14] ), .op(
        n12075) );
  nand2_1 U13607 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][14] ), .op(
        n12074) );
  nand2_1 U13608 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][14] ), .op(
        n12081) );
  nand2_1 U13609 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][14] ), .op(
        n12080) );
  nand2_1 U13610 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][14] ), .op(
        n12079) );
  nand2_1 U13611 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][14] ), .op(
        n12078) );
  inv_1 U13612 ( .ip(n13441), .op(n12880) );
  nor2_1 U13613 ( .ip1(n17765), .ip2(n12836), .op(n12092) );
  nor2_1 U13614 ( .ip1(n12320), .ip2(n12092), .op(n12093) );
  nand2_1 U13615 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][14] ), .op(
        n12096) );
  nand2_1 U13616 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][14] ), .op(
        n12095) );
  nand2_1 U13617 ( .ip1(n12096), .ip2(n12095), .op(n12102) );
  nand2_1 U13618 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][14] ), .op(
        n12100) );
  nand2_1 U13619 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][14] ), .op(
        n12099) );
  nand2_1 U13620 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][14] ), .op(
        n12098) );
  nand2_1 U13621 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][14] ), .op(
        n12097) );
  not_ab_or_c_or_d U13622 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][14] ), .ip3(n12102), .ip4(n12101), .op(n12134) );
  nand2_1 U13623 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][14] ), .op(
        n12106) );
  nand2_1 U13624 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][14] ), .op(
        n12105) );
  nand2_1 U13625 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][14] ), .op(
        n12104) );
  nand2_1 U13626 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][14] ), .op(
        n12103) );
  and4_1 U13627 ( .ip1(n12106), .ip2(n12105), .ip3(n12104), .ip4(n12103), .op(
        n12133) );
  nand2_1 U13628 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][14] ), .op(
        n12110) );
  nand2_1 U13629 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][14] ), .op(
        n12109) );
  nand2_1 U13630 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][14] ), .op(
        n12108) );
  nand2_1 U13631 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][14] ), .op(
        n12107) );
  and4_1 U13632 ( .ip1(n12110), .ip2(n12109), .ip3(n12108), .ip4(n12107), .op(
        n12132) );
  nand2_1 U13633 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][14] ), .op(
        n12114) );
  nand2_1 U13634 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][14] ), .op(
        n12113) );
  nand2_1 U13635 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][14] ), .op(
        n12112) );
  nand2_1 U13636 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][14] ), .op(
        n12111) );
  nand2_1 U13637 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][14] ), .op(
        n12118) );
  nand2_1 U13638 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][14] ), .op(
        n12117) );
  nand2_1 U13639 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][14] ), .op(
        n12116) );
  nand2_1 U13640 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][14] ), .op(
        n12115) );
  nand2_1 U13641 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][14] ), .op(
        n12122) );
  nand2_1 U13642 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][14] ), .op(
        n12121) );
  nand2_1 U13643 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][14] ), .op(
        n12120) );
  nand2_1 U13644 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][14] ), .op(
        n12119) );
  nand2_1 U13645 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][14] ), .op(
        n12126) );
  nand2_1 U13646 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][14] ), .op(
        n12125) );
  nand2_1 U13647 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][14] ), .op(
        n12124) );
  nand2_1 U13648 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][14] ), .op(
        n12123) );
  mux2_1 U13649 ( .ip1(n19330), .ip2(n12135), .s(n13162), .op(n15693) );
  nand2_1 U13650 ( .ip1(n15693), .ip2(n13520), .op(n12137) );
  nand2_1 U13651 ( .ip1(n13521), .ip2(\pipeline/PC_DX [14]), .op(n12136) );
  nand2_1 U13652 ( .ip1(n13636), .ip2(n19432), .op(n13960) );
  nand2_1 U13653 ( .ip1(n13521), .ip2(\pipeline/PC_DX [13]), .op(n12187) );
  nand2_1 U13654 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [13]), .op(n12143) );
  nand2_1 U13655 ( .ip1(\pipeline/alu_out_WB [13]), .ip2(n17895), .op(n12142)
         );
  nand2_1 U13656 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [13]), .op(
        n12141) );
  nand3_1 U13657 ( .ip1(n12143), .ip2(n12142), .ip3(n12141), .op(n19342) );
  nand2_1 U13658 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][13] ), .op(
        n12145) );
  nand2_1 U13659 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][13] ), .op(
        n12144) );
  nand2_1 U13660 ( .ip1(n12145), .ip2(n12144), .op(n12151) );
  nand2_1 U13661 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][13] ), .op(
        n12149) );
  nand2_1 U13662 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][13] ), .op(
        n12148) );
  nand2_1 U13663 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][13] ), .op(
        n12147) );
  nand2_1 U13664 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][13] ), .op(
        n12146) );
  not_ab_or_c_or_d U13665 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][13] ), .ip3(n12151), .ip4(n12150), .op(n12183) );
  nand2_1 U13666 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][13] ), .op(
        n12155) );
  nand2_1 U13667 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][13] ), .op(
        n12154) );
  nand2_1 U13668 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][13] ), .op(
        n12153) );
  nand2_1 U13669 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][13] ), .op(
        n12152) );
  and4_1 U13670 ( .ip1(n12155), .ip2(n12154), .ip3(n12153), .ip4(n12152), .op(
        n12182) );
  nand2_1 U13671 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][13] ), .op(
        n12159) );
  nand2_1 U13672 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][13] ), .op(
        n12158) );
  nand2_1 U13673 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][13] ), .op(
        n12157) );
  nand2_1 U13674 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][13] ), .op(
        n12156) );
  and4_1 U13675 ( .ip1(n12159), .ip2(n12158), .ip3(n12157), .ip4(n12156), .op(
        n12181) );
  nand2_1 U13676 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][13] ), .op(
        n12163) );
  nand2_1 U13677 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][13] ), .op(
        n12162) );
  nand2_1 U13678 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][13] ), .op(
        n12161) );
  nand2_1 U13679 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][13] ), .op(
        n12160) );
  nand2_1 U13680 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][13] ), .op(
        n12167) );
  nand2_1 U13681 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][13] ), .op(
        n12166) );
  nand2_1 U13682 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][13] ), .op(
        n12165) );
  nand2_1 U13683 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][13] ), .op(
        n12164) );
  nand2_1 U13684 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][13] ), .op(
        n12171) );
  nand2_1 U13685 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][13] ), .op(
        n12170) );
  nand2_1 U13686 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][13] ), .op(
        n12169) );
  nand2_1 U13687 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][13] ), .op(
        n12168) );
  nand2_1 U13688 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][13] ), .op(
        n12175) );
  nand2_1 U13689 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][13] ), .op(
        n12174) );
  nand2_1 U13690 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][13] ), .op(
        n12173) );
  nand2_1 U13691 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][13] ), .op(
        n12172) );
  mux2_1 U13692 ( .ip1(n19342), .ip2(n12185), .s(n10200), .op(n20400) );
  nand2_1 U13693 ( .ip1(n20400), .ip2(n13520), .op(n12186) );
  nand2_1 U13694 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][13] ), .op(
        n12189) );
  nand2_1 U13695 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][13] ), .op(
        n12188) );
  nand2_1 U13696 ( .ip1(n12189), .ip2(n12188), .op(n12195) );
  nand2_1 U13697 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][13] ), .op(
        n12193) );
  nand2_1 U13698 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][13] ), .op(
        n12192) );
  nand2_1 U13699 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][13] ), .op(
        n12191) );
  nand2_1 U13700 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][13] ), .op(
        n12190) );
  not_ab_or_c_or_d U13701 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][13] ), .ip3(n12195), .ip4(n12194), .op(n12227) );
  nand2_1 U13702 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][13] ), .op(
        n12199) );
  nand2_1 U13703 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][13] ), .op(
        n12198) );
  nand2_1 U13704 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][13] ), .op(
        n12197) );
  nand2_1 U13705 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][13] ), .op(
        n12196) );
  and4_1 U13706 ( .ip1(n12199), .ip2(n12198), .ip3(n12197), .ip4(n12196), .op(
        n12226) );
  nand2_1 U13707 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][13] ), .op(
        n12203) );
  nand2_1 U13708 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][13] ), .op(
        n12202) );
  nand2_1 U13709 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][13] ), .op(
        n12201) );
  nand2_1 U13710 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][13] ), .op(
        n12200) );
  and4_1 U13711 ( .ip1(n12203), .ip2(n12202), .ip3(n12201), .ip4(n12200), .op(
        n12225) );
  nand2_1 U13712 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][13] ), .op(
        n12207) );
  nand2_1 U13713 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][13] ), .op(
        n12206) );
  nand2_1 U13714 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][13] ), .op(
        n12205) );
  nand2_1 U13715 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][13] ), .op(
        n12204) );
  nand2_1 U13716 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][13] ), .op(
        n12211) );
  nand2_1 U13717 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][13] ), .op(
        n12210) );
  nand2_1 U13718 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][13] ), .op(
        n12209) );
  nand2_1 U13719 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][13] ), .op(
        n12208) );
  nand2_1 U13720 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][13] ), .op(
        n12215) );
  nand2_1 U13721 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][13] ), .op(
        n12214) );
  nand2_1 U13722 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][13] ), .op(
        n12213) );
  nand2_1 U13723 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][13] ), .op(
        n12212) );
  nand2_1 U13724 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][13] ), .op(
        n12219) );
  nand2_1 U13725 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][13] ), .op(
        n12218) );
  nand2_1 U13726 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][13] ), .op(
        n12217) );
  nand2_1 U13727 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][13] ), .op(
        n12216) );
  nor2_1 U13728 ( .ip1(n15352), .ip2(n12836), .op(n12229) );
  nor2_1 U13729 ( .ip1(n12320), .ip2(n12229), .op(n12230) );
  nand2_1 U13730 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [12]), .op(n12234) );
  nand2_1 U13731 ( .ip1(\pipeline/alu_out_WB [12]), .ip2(n17895), .op(n12233)
         );
  nand2_1 U13732 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [12]), .op(
        n12232) );
  nand3_1 U13733 ( .ip1(n12234), .ip2(n12233), .ip3(n12232), .op(n19346) );
  nand2_1 U13734 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][12] ), .op(
        n12236) );
  nand2_1 U13735 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][12] ), .op(
        n12235) );
  nand2_1 U13736 ( .ip1(n12236), .ip2(n12235), .op(n12242) );
  nand2_1 U13737 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][12] ), .op(
        n12240) );
  nand2_1 U13738 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][12] ), .op(
        n12239) );
  nand2_1 U13739 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][12] ), .op(
        n12238) );
  nand2_1 U13740 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][12] ), .op(
        n12237) );
  not_ab_or_c_or_d U13741 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][12] ), .ip3(n12242), .ip4(n12241), .op(n12274) );
  nand2_1 U13742 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][12] ), .op(
        n12246) );
  nand2_1 U13743 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][12] ), .op(
        n12245) );
  nand2_1 U13744 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][12] ), .op(
        n12244) );
  nand2_1 U13745 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][12] ), .op(
        n12243) );
  and4_1 U13746 ( .ip1(n12246), .ip2(n12245), .ip3(n12244), .ip4(n12243), .op(
        n12273) );
  nand2_1 U13747 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][12] ), .op(
        n12250) );
  nand2_1 U13748 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][12] ), .op(
        n12249) );
  nand2_1 U13749 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][12] ), .op(
        n12248) );
  nand2_1 U13750 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][12] ), .op(
        n12247) );
  and4_1 U13751 ( .ip1(n12250), .ip2(n12249), .ip3(n12248), .ip4(n12247), .op(
        n12272) );
  nand2_1 U13752 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][12] ), .op(
        n12254) );
  nand2_1 U13753 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][12] ), .op(
        n12253) );
  nand2_1 U13754 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][12] ), .op(
        n12252) );
  nand2_1 U13755 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][12] ), .op(
        n12251) );
  nand2_1 U13756 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][12] ), .op(
        n12258) );
  nand2_1 U13757 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][12] ), .op(
        n12257) );
  nand2_1 U13758 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][12] ), .op(
        n12256) );
  nand2_1 U13759 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][12] ), .op(
        n12255) );
  nand2_1 U13760 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][12] ), .op(
        n12262) );
  nand2_1 U13761 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][12] ), .op(
        n12261) );
  nand2_1 U13762 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][12] ), .op(
        n12260) );
  nand2_1 U13763 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][12] ), .op(
        n12259) );
  nand2_1 U13764 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][12] ), .op(
        n12266) );
  nand2_1 U13765 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][12] ), .op(
        n12265) );
  nand2_1 U13766 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][12] ), .op(
        n12264) );
  nand2_1 U13767 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][12] ), .op(
        n12263) );
  mux2_1 U13768 ( .ip1(n19346), .ip2(n12275), .s(n10200), .op(n16402) );
  nand2_1 U13769 ( .ip1(n16402), .ip2(n13520), .op(n12277) );
  nand2_1 U13770 ( .ip1(n13521), .ip2(\pipeline/PC_DX [12]), .op(n12276) );
  nand2_1 U13771 ( .ip1(n12277), .ip2(n12276), .op(n13627) );
  nand2_1 U13772 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][12] ), .op(
        n12279) );
  nand2_1 U13773 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][12] ), .op(
        n12278) );
  nand2_1 U13774 ( .ip1(n12279), .ip2(n12278), .op(n12285) );
  nand2_1 U13775 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][12] ), .op(
        n12283) );
  nand2_1 U13776 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][12] ), .op(
        n12282) );
  nand2_1 U13777 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][12] ), .op(
        n12281) );
  nand2_1 U13778 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][12] ), .op(
        n12280) );
  not_ab_or_c_or_d U13779 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][12] ), .ip3(n12285), .ip4(n12284), .op(n12317) );
  nand2_1 U13780 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][12] ), .op(
        n12289) );
  nand2_1 U13781 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][12] ), .op(
        n12288) );
  nand2_1 U13782 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][12] ), .op(
        n12287) );
  nand2_1 U13783 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][12] ), .op(
        n12286) );
  and4_1 U13784 ( .ip1(n12289), .ip2(n12288), .ip3(n12287), .ip4(n12286), .op(
        n12316) );
  nand2_1 U13785 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][12] ), .op(
        n12293) );
  nand2_1 U13786 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][12] ), .op(
        n12292) );
  nand2_1 U13787 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][12] ), .op(
        n12291) );
  nand2_1 U13788 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][12] ), .op(
        n12290) );
  and4_1 U13789 ( .ip1(n12293), .ip2(n12292), .ip3(n12291), .ip4(n12290), .op(
        n12315) );
  nand2_1 U13790 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][12] ), .op(
        n12297) );
  nand2_1 U13791 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][12] ), .op(
        n12296) );
  nand2_1 U13792 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][12] ), .op(
        n12295) );
  nand2_1 U13793 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][12] ), .op(
        n12294) );
  nand2_1 U13794 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][12] ), .op(
        n12301) );
  nand2_1 U13795 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][12] ), .op(
        n12300) );
  nand2_1 U13796 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][12] ), .op(
        n12299) );
  nand2_1 U13797 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][12] ), .op(
        n12298) );
  nand2_1 U13798 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][12] ), .op(
        n12305) );
  nand2_1 U13799 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][12] ), .op(
        n12304) );
  nand2_1 U13800 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][12] ), .op(
        n12303) );
  nand2_1 U13801 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][12] ), .op(
        n12302) );
  nand2_1 U13802 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][12] ), .op(
        n12309) );
  nand2_1 U13803 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][12] ), .op(
        n12308) );
  nand2_1 U13804 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][12] ), .op(
        n12307) );
  nand2_1 U13805 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][12] ), .op(
        n12306) );
  mux2_1 U13806 ( .ip1(n19346), .ip2(n12318), .s(n12683), .op(n22060) );
  nand2_1 U13807 ( .ip1(n22060), .ip2(n10201), .op(n12322) );
  nor2_1 U13808 ( .ip1(n15312), .ip2(n12836), .op(n12319) );
  nor2_1 U13809 ( .ip1(n12320), .ip2(n12319), .op(n12321) );
  nand2_1 U13810 ( .ip1(n12322), .ip2(n12321), .op(n20728) );
  nand2_1 U13811 ( .ip1(n10189), .ip2(n20728), .op(n13626) );
  nor2_1 U13812 ( .ip1(n13678), .ip2(n20222), .op(n12689) );
  or2_1 U13813 ( .ip1(n13626), .ip2(n12689), .op(n12323) );
  nand2_1 U13814 ( .ip1(n13863), .ip2(n12323), .op(n12324) );
  nand2_1 U13815 ( .ip1(n12691), .ip2(n12324), .op(n12325) );
  and2_1 U13816 ( .ip1(n12326), .ip2(n12325), .op(n13833) );
  nand2_1 U13817 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [10]), .op(n12329) );
  nand2_1 U13818 ( .ip1(\pipeline/alu_out_WB [10]), .ip2(n17895), .op(n12328)
         );
  nand2_1 U13819 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [10]), .op(
        n12327) );
  nand3_1 U13820 ( .ip1(n12329), .ip2(n12328), .ip3(n12327), .op(n19396) );
  nand2_1 U13821 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][10] ), .op(
        n12331) );
  nand2_1 U13822 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][10] ), .op(
        n12330) );
  nand2_1 U13823 ( .ip1(n12331), .ip2(n12330), .op(n12337) );
  nand2_1 U13824 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][10] ), .op(
        n12335) );
  nand2_1 U13825 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][10] ), .op(
        n12334) );
  nand2_1 U13826 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][10] ), .op(
        n12333) );
  nand2_1 U13827 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][10] ), .op(
        n12332) );
  not_ab_or_c_or_d U13828 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][10] ), .ip3(n12337), .ip4(n12336), .op(n12369) );
  nand2_1 U13829 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][10] ), .op(
        n12341) );
  nand2_1 U13830 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][10] ), .op(
        n12340) );
  nand2_1 U13831 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][10] ), .op(
        n12339) );
  nand2_1 U13832 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][10] ), .op(
        n12338) );
  and4_1 U13833 ( .ip1(n12341), .ip2(n12340), .ip3(n12339), .ip4(n12338), .op(
        n12368) );
  nand2_1 U13834 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][10] ), .op(
        n12345) );
  nand2_1 U13835 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][10] ), .op(
        n12344) );
  nand2_1 U13836 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][10] ), .op(
        n12343) );
  nand2_1 U13837 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][10] ), .op(
        n12342) );
  and4_1 U13838 ( .ip1(n12345), .ip2(n12344), .ip3(n12343), .ip4(n12342), .op(
        n12367) );
  nand2_1 U13839 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][10] ), .op(
        n12349) );
  nand2_1 U13840 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][10] ), .op(
        n12348) );
  nand2_1 U13841 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][10] ), .op(
        n12347) );
  nand2_1 U13842 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][10] ), .op(
        n12346) );
  nand2_1 U13843 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][10] ), .op(
        n12353) );
  nand2_1 U13844 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][10] ), .op(
        n12352) );
  nand2_1 U13845 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][10] ), .op(
        n12351) );
  nand2_1 U13846 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][10] ), .op(
        n12350) );
  nand2_1 U13847 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][10] ), .op(
        n12357) );
  nand2_1 U13848 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][10] ), .op(
        n12356) );
  nand2_1 U13849 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][10] ), .op(
        n12355) );
  nand2_1 U13850 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][10] ), .op(
        n12354) );
  nand2_1 U13851 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][10] ), .op(
        n12361) );
  nand2_1 U13852 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][10] ), .op(
        n12360) );
  nand2_1 U13853 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][10] ), .op(
        n12359) );
  nand2_1 U13854 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][10] ), .op(
        n12358) );
  mux2_1 U13855 ( .ip1(n19396), .ip2(n12370), .s(n10200), .op(n14601) );
  nand2_1 U13856 ( .ip1(n14601), .ip2(n13520), .op(n12372) );
  nand2_1 U13857 ( .ip1(n13521), .ip2(\pipeline/PC_DX [10]), .op(n12371) );
  nand2_1 U13858 ( .ip1(n12372), .ip2(n12371), .op(n13707) );
  inv_1 U13859 ( .ip(n13707), .op(n13553) );
  nand2_1 U13860 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][10] ), .op(
        n12374) );
  nand2_1 U13861 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][10] ), .op(
        n12373) );
  nand2_1 U13862 ( .ip1(n12374), .ip2(n12373), .op(n12380) );
  nand2_1 U13863 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][10] ), .op(
        n12378) );
  nand2_1 U13864 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][10] ), .op(
        n12377) );
  nand2_1 U13865 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][10] ), .op(
        n12376) );
  nand2_1 U13866 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][10] ), .op(
        n12375) );
  not_ab_or_c_or_d U13867 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][10] ), .ip3(n12380), .ip4(n12379), .op(n12412) );
  nand2_1 U13868 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][10] ), .op(
        n12384) );
  nand2_1 U13869 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][10] ), .op(
        n12383) );
  nand2_1 U13870 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][10] ), .op(
        n12382) );
  nand2_1 U13871 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][10] ), .op(
        n12381) );
  and4_1 U13872 ( .ip1(n12384), .ip2(n12383), .ip3(n12382), .ip4(n12381), .op(
        n12411) );
  nand2_1 U13873 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][10] ), .op(
        n12388) );
  nand2_1 U13874 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][10] ), .op(
        n12387) );
  nand2_1 U13875 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][10] ), .op(
        n12386) );
  nand2_1 U13876 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][10] ), .op(
        n12385) );
  and4_1 U13877 ( .ip1(n12388), .ip2(n12387), .ip3(n12386), .ip4(n12385), .op(
        n12410) );
  nand2_1 U13878 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][10] ), .op(
        n12392) );
  nand2_1 U13879 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][10] ), .op(
        n12391) );
  nand2_1 U13880 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][10] ), .op(
        n12390) );
  nand2_1 U13881 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][10] ), .op(
        n12389) );
  nand2_1 U13882 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][10] ), .op(
        n12396) );
  nand2_1 U13883 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][10] ), .op(
        n12395) );
  nand2_1 U13884 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][10] ), .op(
        n12394) );
  nand2_1 U13885 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][10] ), .op(
        n12393) );
  nand2_1 U13886 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][10] ), .op(
        n12400) );
  nand2_1 U13887 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][10] ), .op(
        n12399) );
  nand2_1 U13888 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][10] ), .op(
        n12398) );
  nand2_1 U13889 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][10] ), .op(
        n12397) );
  nand2_1 U13890 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][10] ), .op(
        n12404) );
  nand2_1 U13891 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][10] ), .op(
        n12403) );
  nand2_1 U13892 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][10] ), .op(
        n12402) );
  nand2_1 U13893 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][10] ), .op(
        n12401) );
  nand2_1 U13894 ( .ip1(n22056), .ip2(n10201), .op(n12415) );
  nand2_1 U13895 ( .ip1(\pipeline/inst_DX [30]), .ip2(n13445), .op(n12414) );
  nor2_1 U13896 ( .ip1(n13553), .ip2(n16972), .op(n13927) );
  nand2_1 U13897 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [11]), .op(n12418) );
  nand2_1 U13898 ( .ip1(\pipeline/alu_out_WB [11]), .ip2(n17895), .op(n12417)
         );
  nand2_1 U13899 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [11]), .op(
        n12416) );
  nand3_1 U13900 ( .ip1(n12418), .ip2(n12417), .ip3(n12416), .op(n19392) );
  nand2_1 U13901 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][11] ), .op(
        n12420) );
  nand2_1 U13902 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][11] ), .op(
        n12419) );
  nand2_1 U13903 ( .ip1(n12420), .ip2(n12419), .op(n12426) );
  nand2_1 U13904 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][11] ), .op(
        n12424) );
  nand2_1 U13905 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][11] ), .op(
        n12423) );
  nand2_1 U13906 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][11] ), .op(
        n12422) );
  nand2_1 U13907 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][11] ), .op(
        n12421) );
  not_ab_or_c_or_d U13908 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][11] ), .ip3(n12426), .ip4(n12425), .op(n12458) );
  nand2_1 U13909 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][11] ), .op(
        n12430) );
  nand2_1 U13910 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][11] ), .op(
        n12429) );
  nand2_1 U13911 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][11] ), .op(
        n12428) );
  nand2_1 U13912 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][11] ), .op(
        n12427) );
  and4_1 U13913 ( .ip1(n12430), .ip2(n12429), .ip3(n12428), .ip4(n12427), .op(
        n12457) );
  nand2_1 U13914 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][11] ), .op(
        n12434) );
  nand2_1 U13915 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][11] ), .op(
        n12433) );
  nand2_1 U13916 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][11] ), .op(
        n12432) );
  nand2_1 U13917 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][11] ), .op(
        n12431) );
  and4_1 U13918 ( .ip1(n12434), .ip2(n12433), .ip3(n12432), .ip4(n12431), .op(
        n12456) );
  nand2_1 U13919 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][11] ), .op(
        n12438) );
  nand2_1 U13920 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][11] ), .op(
        n12437) );
  nand2_1 U13921 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][11] ), .op(
        n12436) );
  nand2_1 U13922 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][11] ), .op(
        n12435) );
  nand2_1 U13923 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][11] ), .op(
        n12442) );
  nand2_1 U13924 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][11] ), .op(
        n12441) );
  nand2_1 U13925 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][11] ), .op(
        n12440) );
  nand2_1 U13926 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][11] ), .op(
        n12439) );
  nand2_1 U13927 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][11] ), .op(
        n12446) );
  nand2_1 U13928 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][11] ), .op(
        n12445) );
  nand2_1 U13929 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][11] ), .op(
        n12444) );
  nand2_1 U13930 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][11] ), .op(
        n12443) );
  nand2_1 U13931 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][11] ), .op(
        n12450) );
  nand2_1 U13932 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][11] ), .op(
        n12449) );
  nand2_1 U13933 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][11] ), .op(
        n12448) );
  nand2_1 U13934 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][11] ), .op(
        n12447) );
  mux2_1 U13935 ( .ip1(n19392), .ip2(n12459), .s(n10200), .op(n16226) );
  nand2_1 U13936 ( .ip1(n16226), .ip2(n13520), .op(n12461) );
  nand2_1 U13937 ( .ip1(n13521), .ip2(\pipeline/PC_DX [11]), .op(n12460) );
  nand2_1 U13938 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][11] ), .op(
        n12463) );
  nand2_1 U13939 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][11] ), .op(
        n12462) );
  nand2_1 U13940 ( .ip1(n12463), .ip2(n12462), .op(n12469) );
  nand2_1 U13941 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][11] ), .op(
        n12467) );
  nand2_1 U13942 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][11] ), .op(
        n12466) );
  nand2_1 U13943 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][11] ), .op(
        n12465) );
  nand2_1 U13944 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][11] ), .op(
        n12464) );
  not_ab_or_c_or_d U13945 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][11] ), .ip3(n12469), .ip4(n12468), .op(n12501) );
  nand2_1 U13946 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][11] ), .op(
        n12473) );
  nand2_1 U13947 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][11] ), .op(
        n12472) );
  nand2_1 U13948 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][11] ), .op(
        n12471) );
  nand2_1 U13949 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][11] ), .op(
        n12470) );
  and4_1 U13950 ( .ip1(n12473), .ip2(n12472), .ip3(n12471), .ip4(n12470), .op(
        n12500) );
  nand2_1 U13951 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][11] ), .op(
        n12477) );
  nand2_1 U13952 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][11] ), .op(
        n12476) );
  nand2_1 U13953 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][11] ), .op(
        n12475) );
  nand2_1 U13954 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][11] ), .op(
        n12474) );
  and4_1 U13955 ( .ip1(n12477), .ip2(n12476), .ip3(n12475), .ip4(n12474), .op(
        n12499) );
  nand2_1 U13956 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][11] ), .op(
        n12481) );
  nand2_1 U13957 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][11] ), .op(
        n12480) );
  nand2_1 U13958 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][11] ), .op(
        n12479) );
  nand2_1 U13959 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][11] ), .op(
        n12478) );
  nand2_1 U13960 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][11] ), .op(
        n12485) );
  nand2_1 U13961 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][11] ), .op(
        n12484) );
  nand2_1 U13962 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][11] ), .op(
        n12483) );
  nand2_1 U13963 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][11] ), .op(
        n12482) );
  nand2_1 U13964 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][11] ), .op(
        n12489) );
  nand2_1 U13965 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][11] ), .op(
        n12488) );
  nand2_1 U13966 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][11] ), .op(
        n12487) );
  nand2_1 U13967 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][11] ), .op(
        n12486) );
  nand2_1 U13968 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][11] ), .op(
        n12493) );
  nand2_1 U13969 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][11] ), .op(
        n12492) );
  nand2_1 U13970 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][11] ), .op(
        n12491) );
  nand2_1 U13971 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][11] ), .op(
        n12490) );
  mux2_1 U13972 ( .ip1(n19392), .ip2(n12502), .s(n12683), .op(n22058) );
  nand2_1 U13973 ( .ip1(n22058), .ip2(n10201), .op(n12504) );
  nor2_1 U13974 ( .ip1(n13552), .ip2(n16690), .op(n13554) );
  nor2_1 U13975 ( .ip1(n13927), .ip2(n13554), .op(n13559) );
  nand2_1 U13976 ( .ip1(\pipeline/regfile/data[8][8] ), .ip2(n13448), .op(
        n12506) );
  nand2_1 U13977 ( .ip1(\pipeline/regfile/data[10][8] ), .ip2(n13449), .op(
        n12505) );
  nand2_1 U13978 ( .ip1(n12506), .ip2(n12505), .op(n12512) );
  nand2_1 U13979 ( .ip1(\pipeline/regfile/data[21][8] ), .ip2(n13452), .op(
        n12510) );
  nand2_1 U13980 ( .ip1(\pipeline/regfile/data[17][8] ), .ip2(n13453), .op(
        n12509) );
  nand2_1 U13981 ( .ip1(\pipeline/regfile/data[7][8] ), .ip2(n13454), .op(
        n12508) );
  nand2_1 U13982 ( .ip1(\pipeline/regfile/data[1][8] ), .ip2(n13455), .op(
        n12507) );
  not_ab_or_c_or_d U13983 ( .ip1(\pipeline/regfile/data[28][8] ), .ip2(n13462), 
        .ip3(n12512), .ip4(n12511), .op(n12544) );
  nand2_1 U13984 ( .ip1(\pipeline/regfile/data[27][8] ), .ip2(n13463), .op(
        n12516) );
  nand2_1 U13985 ( .ip1(\pipeline/regfile/data[9][8] ), .ip2(n13464), .op(
        n12515) );
  nand2_1 U13986 ( .ip1(\pipeline/regfile/data[2][8] ), .ip2(n13465), .op(
        n12514) );
  nand2_1 U13987 ( .ip1(\pipeline/regfile/data[26][8] ), .ip2(n13466), .op(
        n12513) );
  and4_1 U13988 ( .ip1(n12516), .ip2(n12515), .ip3(n12514), .ip4(n12513), .op(
        n12543) );
  nand2_1 U13989 ( .ip1(\pipeline/regfile/data[16][8] ), .ip2(n13471), .op(
        n12520) );
  nand2_1 U13990 ( .ip1(\pipeline/regfile/data[4][8] ), .ip2(n13472), .op(
        n12519) );
  nand2_1 U13991 ( .ip1(\pipeline/regfile/data[24][8] ), .ip2(n13473), .op(
        n12518) );
  nand2_1 U13992 ( .ip1(\pipeline/regfile/data[20][8] ), .ip2(n13474), .op(
        n12517) );
  and4_1 U13993 ( .ip1(n12520), .ip2(n12519), .ip3(n12518), .ip4(n12517), .op(
        n12542) );
  nand2_1 U13994 ( .ip1(\pipeline/regfile/data[25][8] ), .ip2(n13479), .op(
        n12524) );
  nand2_1 U13995 ( .ip1(\pipeline/regfile/data[3][8] ), .ip2(n13480), .op(
        n12523) );
  nand2_1 U13996 ( .ip1(\pipeline/regfile/data[6][8] ), .ip2(n13481), .op(
        n12522) );
  nand2_1 U13997 ( .ip1(\pipeline/regfile/data[5][8] ), .ip2(n13482), .op(
        n12521) );
  nand2_1 U13998 ( .ip1(\pipeline/regfile/data[18][8] ), .ip2(n13487), .op(
        n12528) );
  nand2_1 U13999 ( .ip1(\pipeline/regfile/data[23][8] ), .ip2(n13488), .op(
        n12527) );
  nand2_1 U14000 ( .ip1(\pipeline/regfile/data[11][8] ), .ip2(n13489), .op(
        n12526) );
  nand2_1 U14001 ( .ip1(\pipeline/regfile/data[19][8] ), .ip2(n13490), .op(
        n12525) );
  nand2_1 U14002 ( .ip1(\pipeline/regfile/data[29][8] ), .ip2(n13495), .op(
        n12532) );
  nand2_1 U14003 ( .ip1(\pipeline/regfile/data[22][8] ), .ip2(n13496), .op(
        n12531) );
  nand2_1 U14004 ( .ip1(\pipeline/regfile/data[15][8] ), .ip2(n13497), .op(
        n12530) );
  nand2_1 U14005 ( .ip1(\pipeline/regfile/data[31][8] ), .ip2(n13498), .op(
        n12529) );
  nand2_1 U14006 ( .ip1(\pipeline/regfile/data[14][8] ), .ip2(n13503), .op(
        n12536) );
  nand2_1 U14007 ( .ip1(\pipeline/regfile/data[13][8] ), .ip2(n13504), .op(
        n12535) );
  nand2_1 U14008 ( .ip1(\pipeline/regfile/data[30][8] ), .ip2(n13505), .op(
        n12534) );
  nand2_1 U14009 ( .ip1(\pipeline/regfile/data[12][8] ), .ip2(n13506), .op(
        n12533) );
  and4_1 U14010 ( .ip1(n12544), .ip2(n12543), .ip3(n12542), .ip4(n12541), .op(
        n12545) );
  nand2_1 U14011 ( .ip1(n14057), .ip2(n12545), .op(n14122) );
  nand2_1 U14012 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [8]), .op(n12548)
         );
  nand2_1 U14013 ( .ip1(\pipeline/alu_out_WB [8]), .ip2(n17895), .op(n12547)
         );
  nand2_1 U14014 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [8]), .op(
        n12546) );
  nand3_1 U14015 ( .ip1(n12548), .ip2(n12547), .ip3(n12546), .op(n12592) );
  inv_1 U14016 ( .ip(n12592), .op(n19405) );
  nand2_1 U14017 ( .ip1(n12549), .ip2(n19405), .op(n14121) );
  nand3_1 U14018 ( .ip1(n14122), .ip2(n13520), .ip3(n14121), .op(n12551) );
  nand2_1 U14019 ( .ip1(n13521), .ip2(\pipeline/PC_DX [8]), .op(n12550) );
  nand2_1 U14020 ( .ip1(n12551), .ip2(n12550), .op(n13698) );
  nand2_1 U14021 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][8] ), .op(
        n12553) );
  nand2_1 U14022 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][8] ), .op(
        n12552) );
  nand2_1 U14023 ( .ip1(n12553), .ip2(n12552), .op(n12559) );
  nand2_1 U14024 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][8] ), .op(
        n12557) );
  nand2_1 U14025 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][8] ), .op(
        n12556) );
  nand2_1 U14026 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][8] ), .op(
        n12555) );
  nand2_1 U14027 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][8] ), .op(
        n12554) );
  not_ab_or_c_or_d U14028 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][8] ), 
        .ip3(n12559), .ip4(n12558), .op(n12591) );
  nand2_1 U14029 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][8] ), .op(
        n12563) );
  nand2_1 U14030 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][8] ), .op(
        n12562) );
  nand2_1 U14031 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][8] ), .op(
        n12561) );
  nand2_1 U14032 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][8] ), .op(
        n12560) );
  and4_1 U14033 ( .ip1(n12563), .ip2(n12562), .ip3(n12561), .ip4(n12560), .op(
        n12590) );
  nand2_1 U14034 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][8] ), .op(
        n12567) );
  nand2_1 U14035 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][8] ), .op(
        n12566) );
  nand2_1 U14036 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][8] ), .op(
        n12565) );
  nand2_1 U14037 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][8] ), .op(
        n12564) );
  and4_1 U14038 ( .ip1(n12567), .ip2(n12566), .ip3(n12565), .ip4(n12564), .op(
        n12589) );
  nand2_1 U14039 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][8] ), .op(
        n12571) );
  nand2_1 U14040 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][8] ), .op(
        n12570) );
  nand2_1 U14041 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][8] ), .op(
        n12569) );
  nand2_1 U14042 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][8] ), .op(
        n12568) );
  nand2_1 U14043 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][8] ), .op(
        n12575) );
  nand2_1 U14044 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][8] ), .op(
        n12574) );
  nand2_1 U14045 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][8] ), .op(
        n12573) );
  nand2_1 U14046 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][8] ), .op(
        n12572) );
  nand2_1 U14047 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][8] ), .op(
        n12579) );
  nand2_1 U14048 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][8] ), .op(
        n12578) );
  nand2_1 U14049 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][8] ), .op(
        n12577) );
  nand2_1 U14050 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][8] ), .op(
        n12576) );
  nand2_1 U14051 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][8] ), .op(
        n12583) );
  nand2_1 U14052 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][8] ), .op(
        n12582) );
  nand2_1 U14053 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][8] ), .op(
        n12581) );
  nand2_1 U14054 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][8] ), .op(
        n12580) );
  mux2_1 U14055 ( .ip1(n12593), .ip2(n12592), .s(n12880), .op(n22052) );
  nand2_1 U14056 ( .ip1(\pipeline/inst_DX [28]), .ip2(n13445), .op(n12594) );
  nor2_1 U14057 ( .ip1(n16811), .ip2(n12596), .op(n12687) );
  nand2_1 U14058 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [9]), .op(n12599)
         );
  nand2_1 U14059 ( .ip1(\pipeline/alu_out_WB [9]), .ip2(n17895), .op(n12598)
         );
  nand2_1 U14060 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [9]), .op(
        n12597) );
  nand3_1 U14061 ( .ip1(n12599), .ip2(n12598), .ip3(n12597), .op(n18423) );
  nand2_1 U14062 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][9] ), .op(
        n12601) );
  nand2_1 U14063 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][9] ), .op(
        n12600) );
  nand2_1 U14064 ( .ip1(n12601), .ip2(n12600), .op(n12607) );
  nand2_1 U14065 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][9] ), .op(
        n12605) );
  nand2_1 U14066 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][9] ), .op(
        n12604) );
  nand2_1 U14067 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][9] ), .op(
        n12603) );
  nand2_1 U14068 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][9] ), .op(
        n12602) );
  not_ab_or_c_or_d U14069 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][9] ), 
        .ip3(n12607), .ip4(n12606), .op(n12639) );
  nand2_1 U14070 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][9] ), .op(
        n12611) );
  nand2_1 U14071 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][9] ), .op(
        n12610) );
  nand2_1 U14072 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][9] ), .op(
        n12609) );
  nand2_1 U14073 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][9] ), .op(
        n12608) );
  and4_1 U14074 ( .ip1(n12611), .ip2(n12610), .ip3(n12609), .ip4(n12608), .op(
        n12638) );
  nand2_1 U14075 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][9] ), .op(
        n12615) );
  nand2_1 U14076 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][9] ), .op(
        n12614) );
  nand2_1 U14077 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][9] ), .op(
        n12613) );
  nand2_1 U14078 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][9] ), .op(
        n12612) );
  and4_1 U14079 ( .ip1(n12615), .ip2(n12614), .ip3(n12613), .ip4(n12612), .op(
        n12637) );
  nand2_1 U14080 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][9] ), .op(
        n12619) );
  nand2_1 U14081 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][9] ), .op(
        n12618) );
  nand2_1 U14082 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][9] ), .op(
        n12617) );
  nand2_1 U14083 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][9] ), .op(
        n12616) );
  nand2_1 U14084 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][9] ), .op(
        n12623) );
  nand2_1 U14085 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][9] ), .op(
        n12622) );
  nand2_1 U14086 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][9] ), .op(
        n12621) );
  nand2_1 U14087 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][9] ), .op(
        n12620) );
  nand2_1 U14088 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][9] ), .op(
        n12627) );
  nand2_1 U14089 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][9] ), .op(
        n12626) );
  nand2_1 U14090 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][9] ), .op(
        n12625) );
  nand2_1 U14091 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][9] ), .op(
        n12624) );
  nand2_1 U14092 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][9] ), .op(
        n12631) );
  nand2_1 U14093 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][9] ), .op(
        n12630) );
  nand2_1 U14094 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][9] ), .op(
        n12629) );
  nand2_1 U14095 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][9] ), .op(
        n12628) );
  mux2_1 U14096 ( .ip1(n18423), .ip2(n12640), .s(n14057), .op(n15896) );
  nand2_1 U14097 ( .ip1(n15896), .ip2(n13520), .op(n12642) );
  nand2_1 U14098 ( .ip1(n13521), .ip2(\pipeline/PC_DX [9]), .op(n12641) );
  nand2_1 U14099 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][9] ), .op(
        n12644) );
  nand2_1 U14100 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][9] ), .op(
        n12643) );
  nand2_1 U14101 ( .ip1(n12644), .ip2(n12643), .op(n12650) );
  nand2_1 U14102 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][9] ), .op(
        n12648) );
  nand2_1 U14103 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][9] ), .op(
        n12647) );
  nand2_1 U14104 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][9] ), .op(
        n12646) );
  nand2_1 U14105 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][9] ), .op(
        n12645) );
  not_ab_or_c_or_d U14106 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][9] ), 
        .ip3(n12650), .ip4(n12649), .op(n12682) );
  nand2_1 U14107 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][9] ), .op(
        n12654) );
  nand2_1 U14108 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][9] ), .op(
        n12653) );
  nand2_1 U14109 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][9] ), .op(
        n12652) );
  nand2_1 U14110 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][9] ), .op(
        n12651) );
  and4_1 U14111 ( .ip1(n12654), .ip2(n12653), .ip3(n12652), .ip4(n12651), .op(
        n12681) );
  nand2_1 U14112 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][9] ), .op(
        n12658) );
  nand2_1 U14113 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][9] ), .op(
        n12657) );
  nand2_1 U14114 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][9] ), .op(
        n12656) );
  nand2_1 U14115 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][9] ), .op(
        n12655) );
  and4_1 U14116 ( .ip1(n12658), .ip2(n12657), .ip3(n12656), .ip4(n12655), .op(
        n12680) );
  nand2_1 U14117 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][9] ), .op(
        n12662) );
  nand2_1 U14118 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][9] ), .op(
        n12661) );
  nand2_1 U14119 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][9] ), .op(
        n12660) );
  nand2_1 U14120 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][9] ), .op(
        n12659) );
  nand2_1 U14121 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][9] ), .op(
        n12666) );
  nand2_1 U14122 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][9] ), .op(
        n12665) );
  nand2_1 U14123 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][9] ), .op(
        n12664) );
  nand2_1 U14124 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][9] ), .op(
        n12663) );
  nand2_1 U14125 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][9] ), .op(
        n12670) );
  nand2_1 U14126 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][9] ), .op(
        n12669) );
  nand2_1 U14127 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][9] ), .op(
        n12668) );
  nand2_1 U14128 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][9] ), .op(
        n12667) );
  nand2_1 U14129 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][9] ), .op(
        n12674) );
  nand2_1 U14130 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][9] ), .op(
        n12673) );
  nand2_1 U14131 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][9] ), .op(
        n12672) );
  nand2_1 U14132 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][9] ), .op(
        n12671) );
  nand2_1 U14133 ( .ip1(n22054), .ip2(n10201), .op(n12686) );
  nand2_1 U14134 ( .ip1(n13445), .ip2(\pipeline/inst_DX [29]), .op(n12685) );
  nor2_1 U14135 ( .ip1(n12687), .ip2(n13925), .op(n12688) );
  nand2_1 U14136 ( .ip1(n13559), .ip2(n12688), .op(n12693) );
  nor2_1 U14137 ( .ip1(n10189), .ip2(n20728), .op(n12690) );
  nor2_1 U14138 ( .ip1(n12690), .ip2(n12689), .op(n12692) );
  nor2_1 U14139 ( .ip1(n12693), .ip2(n13832), .op(n13551) );
  nand2_1 U14140 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [5]), .op(n12696)
         );
  nand2_1 U14141 ( .ip1(\pipeline/alu_out_WB [5]), .ip2(n17895), .op(n12695)
         );
  nand2_1 U14142 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [5]), .op(
        n12694) );
  nand3_1 U14143 ( .ip1(n12696), .ip2(n12695), .ip3(n12694), .op(n17978) );
  or2_1 U14144 ( .ip1(n12742), .ip2(n13364), .op(n12739) );
  nand2_1 U14145 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][5] ), .op(
        n12698) );
  nand2_1 U14146 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][5] ), .op(
        n12697) );
  nand2_1 U14147 ( .ip1(n12698), .ip2(n12697), .op(n12704) );
  nand2_1 U14148 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][5] ), .op(
        n12702) );
  nand2_1 U14149 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][5] ), .op(
        n12701) );
  nand2_1 U14150 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][5] ), .op(
        n12700) );
  nand2_1 U14151 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][5] ), .op(
        n12699) );
  not_ab_or_c_or_d U14152 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][5] ), 
        .ip3(n12704), .ip4(n12703), .op(n12736) );
  nand2_1 U14153 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][5] ), .op(
        n12708) );
  nand2_1 U14154 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][5] ), .op(
        n12707) );
  nand2_1 U14155 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][5] ), .op(
        n12706) );
  nand2_1 U14156 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][5] ), .op(
        n12705) );
  and4_1 U14157 ( .ip1(n12708), .ip2(n12707), .ip3(n12706), .ip4(n12705), .op(
        n12735) );
  nand2_1 U14158 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][5] ), .op(
        n12712) );
  nand2_1 U14159 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][5] ), .op(
        n12711) );
  nand2_1 U14160 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][5] ), .op(
        n12710) );
  nand2_1 U14161 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][5] ), .op(
        n12709) );
  and4_1 U14162 ( .ip1(n12712), .ip2(n12711), .ip3(n12710), .ip4(n12709), .op(
        n12734) );
  nand2_1 U14163 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][5] ), .op(
        n12716) );
  nand2_1 U14164 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][5] ), .op(
        n12715) );
  nand2_1 U14165 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][5] ), .op(
        n12714) );
  nand2_1 U14166 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][5] ), .op(
        n12713) );
  nand2_1 U14167 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][5] ), .op(
        n12720) );
  nand2_1 U14168 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][5] ), .op(
        n12719) );
  nand2_1 U14169 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][5] ), .op(
        n12718) );
  nand2_1 U14170 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][5] ), .op(
        n12717) );
  nand2_1 U14171 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][5] ), .op(
        n12724) );
  nand2_1 U14172 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][5] ), .op(
        n12723) );
  nand2_1 U14173 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][5] ), .op(
        n12722) );
  nand2_1 U14174 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][5] ), .op(
        n12721) );
  nand2_1 U14175 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][5] ), .op(
        n12728) );
  nand2_1 U14176 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][5] ), .op(
        n12727) );
  nand2_1 U14177 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][5] ), .op(
        n12726) );
  nand2_1 U14178 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][5] ), .op(
        n12725) );
  nand2_1 U14179 ( .ip1(n12737), .ip2(n14057), .op(n12738) );
  nand2_1 U14180 ( .ip1(n12739), .ip2(n12738), .op(n20476) );
  nand2_1 U14181 ( .ip1(n20476), .ip2(n13520), .op(n12741) );
  nand2_1 U14182 ( .ip1(n13521), .ip2(\pipeline/PC_DX [5]), .op(n12740) );
  nand2_1 U14183 ( .ip1(\pipeline/inst_DX [25]), .ip2(n13445), .op(n12787) );
  inv_1 U14184 ( .ip(n17978), .op(n12742) );
  or2_1 U14185 ( .ip1(n12742), .ip2(n13441), .op(n12785) );
  nand2_1 U14186 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][5] ), .op(
        n12744) );
  nand2_1 U14187 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][5] ), .op(
        n12743) );
  nand2_1 U14188 ( .ip1(n12744), .ip2(n12743), .op(n12750) );
  nand2_1 U14189 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][5] ), .op(
        n12748) );
  nand2_1 U14190 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][5] ), .op(
        n12747) );
  nand2_1 U14191 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][5] ), .op(
        n12746) );
  nand2_1 U14192 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][5] ), .op(
        n12745) );
  not_ab_or_c_or_d U14193 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][5] ), 
        .ip3(n12750), .ip4(n12749), .op(n12782) );
  nand2_1 U14194 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][5] ), .op(
        n12754) );
  nand2_1 U14195 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][5] ), .op(
        n12753) );
  nand2_1 U14196 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][5] ), .op(
        n12752) );
  nand2_1 U14197 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][5] ), .op(
        n12751) );
  and4_1 U14198 ( .ip1(n12754), .ip2(n12753), .ip3(n12752), .ip4(n12751), .op(
        n12781) );
  nand2_1 U14199 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][5] ), .op(
        n12758) );
  nand2_1 U14200 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][5] ), .op(
        n12757) );
  nand2_1 U14201 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][5] ), .op(
        n12756) );
  nand2_1 U14202 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][5] ), .op(
        n12755) );
  and4_1 U14203 ( .ip1(n12758), .ip2(n12757), .ip3(n12756), .ip4(n12755), .op(
        n12780) );
  nand2_1 U14204 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][5] ), .op(
        n12762) );
  nand2_1 U14205 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][5] ), .op(
        n12761) );
  nand2_1 U14206 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][5] ), .op(
        n12760) );
  nand2_1 U14207 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][5] ), .op(
        n12759) );
  nand2_1 U14208 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][5] ), .op(
        n12766) );
  nand2_1 U14209 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][5] ), .op(
        n12765) );
  nand2_1 U14210 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][5] ), .op(
        n12764) );
  nand2_1 U14211 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][5] ), .op(
        n12763) );
  nand2_1 U14212 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][5] ), .op(
        n12770) );
  nand2_1 U14213 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][5] ), .op(
        n12769) );
  nand2_1 U14214 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][5] ), .op(
        n12768) );
  nand2_1 U14215 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][5] ), .op(
        n12767) );
  nand2_1 U14216 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][5] ), .op(
        n12774) );
  nand2_1 U14217 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][5] ), .op(
        n12773) );
  nand2_1 U14218 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][5] ), .op(
        n12772) );
  nand2_1 U14219 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][5] ), .op(
        n12771) );
  nand2_1 U14220 ( .ip1(n12783), .ip2(n12683), .op(n12784) );
  nand2_1 U14221 ( .ip1(n12785), .ip2(n12784), .op(n17370) );
  nand2_1 U14222 ( .ip1(n16445), .ip2(n10194), .op(n12788) );
  inv_1 U14223 ( .ip(n12788), .op(n13541) );
  nand2_1 U14224 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [4]), .op(n12791)
         );
  nand2_1 U14225 ( .ip1(\pipeline/alu_out_WB [4]), .ip2(n17895), .op(n12790)
         );
  nand2_1 U14226 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [4]), .op(
        n12789) );
  nand3_1 U14227 ( .ip1(n12791), .ip2(n12790), .ip3(n12789), .op(n17931) );
  nand2_1 U14228 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][4] ), .op(
        n12793) );
  nand2_1 U14229 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][4] ), .op(
        n12792) );
  nand2_1 U14230 ( .ip1(n12793), .ip2(n12792), .op(n12799) );
  nand2_1 U14231 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][4] ), .op(
        n12797) );
  nand2_1 U14232 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][4] ), .op(
        n12796) );
  nand2_1 U14233 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][4] ), .op(
        n12795) );
  nand2_1 U14234 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][4] ), .op(
        n12794) );
  not_ab_or_c_or_d U14235 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][4] ), 
        .ip3(n12799), .ip4(n12798), .op(n12831) );
  nand2_1 U14236 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][4] ), .op(
        n12803) );
  nand2_1 U14237 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][4] ), .op(
        n12802) );
  nand2_1 U14238 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][4] ), .op(
        n12801) );
  nand2_1 U14239 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][4] ), .op(
        n12800) );
  and4_1 U14240 ( .ip1(n12803), .ip2(n12802), .ip3(n12801), .ip4(n12800), .op(
        n12830) );
  nand2_1 U14241 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][4] ), .op(
        n12807) );
  nand2_1 U14242 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][4] ), .op(
        n12806) );
  nand2_1 U14243 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][4] ), .op(
        n12805) );
  nand2_1 U14244 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][4] ), .op(
        n12804) );
  and4_1 U14245 ( .ip1(n12807), .ip2(n12806), .ip3(n12805), .ip4(n12804), .op(
        n12829) );
  nand2_1 U14246 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][4] ), .op(
        n12811) );
  nand2_1 U14247 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][4] ), .op(
        n12810) );
  nand2_1 U14248 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][4] ), .op(
        n12809) );
  nand2_1 U14249 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][4] ), .op(
        n12808) );
  nand2_1 U14250 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][4] ), .op(
        n12815) );
  nand2_1 U14251 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][4] ), .op(
        n12814) );
  nand2_1 U14252 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][4] ), .op(
        n12813) );
  nand2_1 U14253 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][4] ), .op(
        n12812) );
  nand2_1 U14254 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][4] ), .op(
        n12819) );
  nand2_1 U14255 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][4] ), .op(
        n12818) );
  nand2_1 U14256 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][4] ), .op(
        n12817) );
  nand2_1 U14257 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][4] ), .op(
        n12816) );
  nand2_1 U14258 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][4] ), .op(
        n12823) );
  nand2_1 U14259 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][4] ), .op(
        n12822) );
  nand2_1 U14260 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][4] ), .op(
        n12821) );
  nand2_1 U14261 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][4] ), .op(
        n12820) );
  mux2_1 U14262 ( .ip1(n17931), .ip2(n12832), .s(n10200), .op(n17939) );
  nand2_1 U14263 ( .ip1(n17939), .ip2(n13520), .op(n12834) );
  nand2_1 U14264 ( .ip1(n13521), .ip2(\pipeline/PC_DX [4]), .op(n12833) );
  inv_1 U14265 ( .ip(\pipeline/inst_DX [11]), .op(n12835) );
  nor2_1 U14266 ( .ip1(n13443), .ip2(n12835), .op(n12839) );
  nand3_1 U14267 ( .ip1(n13443), .ip2(n13220), .ip3(n12836), .op(n13318) );
  nor2_1 U14268 ( .ip1(n12837), .ip2(n13318), .op(n12838) );
  nor2_1 U14269 ( .ip1(n12839), .ip2(n12838), .op(n12882) );
  nand2_1 U14270 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][4] ), .op(
        n12841) );
  nand2_1 U14271 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][4] ), .op(
        n12840) );
  nand2_1 U14272 ( .ip1(n12841), .ip2(n12840), .op(n12847) );
  nand2_1 U14273 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][4] ), .op(
        n12845) );
  nand2_1 U14274 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][4] ), .op(
        n12844) );
  nand2_1 U14275 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][4] ), .op(
        n12843) );
  nand2_1 U14276 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][4] ), .op(
        n12842) );
  not_ab_or_c_or_d U14277 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][4] ), 
        .ip3(n12847), .ip4(n12846), .op(n12879) );
  nand2_1 U14278 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][4] ), .op(
        n12851) );
  nand2_1 U14279 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][4] ), .op(
        n12850) );
  nand2_1 U14280 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][4] ), .op(
        n12849) );
  nand2_1 U14281 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][4] ), .op(
        n12848) );
  and4_1 U14282 ( .ip1(n12851), .ip2(n12850), .ip3(n12849), .ip4(n12848), .op(
        n12878) );
  nand2_1 U14283 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][4] ), .op(
        n12855) );
  nand2_1 U14284 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][4] ), .op(
        n12854) );
  nand2_1 U14285 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][4] ), .op(
        n12853) );
  nand2_1 U14286 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][4] ), .op(
        n12852) );
  and4_1 U14287 ( .ip1(n12855), .ip2(n12854), .ip3(n12853), .ip4(n12852), .op(
        n12877) );
  nand2_1 U14288 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][4] ), .op(
        n12859) );
  nand2_1 U14289 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][4] ), .op(
        n12858) );
  nand2_1 U14290 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][4] ), .op(
        n12857) );
  nand2_1 U14291 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][4] ), .op(
        n12856) );
  nand2_1 U14292 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][4] ), .op(
        n12863) );
  nand2_1 U14293 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][4] ), .op(
        n12862) );
  nand2_1 U14294 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][4] ), .op(
        n12861) );
  nand2_1 U14295 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][4] ), .op(
        n12860) );
  nand2_1 U14296 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][4] ), .op(
        n12867) );
  nand2_1 U14297 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][4] ), .op(
        n12866) );
  nand2_1 U14298 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][4] ), .op(
        n12865) );
  nand2_1 U14299 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][4] ), .op(
        n12864) );
  nand2_1 U14300 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][4] ), .op(
        n12871) );
  nand2_1 U14301 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][4] ), .op(
        n12870) );
  nand2_1 U14302 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][4] ), .op(
        n12869) );
  nand2_1 U14303 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][4] ), .op(
        n12868) );
  nor2_1 U14304 ( .ip1(n13540), .ip2(n17199), .op(n13913) );
  nor2_1 U14305 ( .ip1(n13541), .ip2(n13913), .op(n13068) );
  nand2_1 U14306 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [6]), .op(n12888)
         );
  nand2_1 U14307 ( .ip1(\pipeline/alu_out_WB [6]), .ip2(n17895), .op(n12887)
         );
  nand2_1 U14308 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [6]), .op(
        n12886) );
  nand3_1 U14309 ( .ip1(n12888), .ip2(n12887), .ip3(n12886), .op(n18007) );
  nand2_1 U14310 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][6] ), .op(
        n12890) );
  nand2_1 U14311 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][6] ), .op(
        n12889) );
  nand2_1 U14312 ( .ip1(n12890), .ip2(n12889), .op(n12896) );
  nand2_1 U14313 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][6] ), .op(
        n12894) );
  nand2_1 U14314 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][6] ), .op(
        n12893) );
  nand2_1 U14315 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][6] ), .op(
        n12892) );
  nand2_1 U14316 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][6] ), .op(
        n12891) );
  not_ab_or_c_or_d U14317 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][6] ), 
        .ip3(n12896), .ip4(n12895), .op(n12928) );
  nand2_1 U14318 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][6] ), .op(
        n12900) );
  nand2_1 U14319 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][6] ), .op(
        n12899) );
  nand2_1 U14320 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][6] ), .op(
        n12898) );
  nand2_1 U14321 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][6] ), .op(
        n12897) );
  and4_1 U14322 ( .ip1(n12900), .ip2(n12899), .ip3(n12898), .ip4(n12897), .op(
        n12927) );
  nand2_1 U14323 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][6] ), .op(
        n12904) );
  nand2_1 U14324 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][6] ), .op(
        n12903) );
  nand2_1 U14325 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][6] ), .op(
        n12902) );
  nand2_1 U14326 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][6] ), .op(
        n12901) );
  and4_1 U14327 ( .ip1(n12904), .ip2(n12903), .ip3(n12902), .ip4(n12901), .op(
        n12926) );
  nand2_1 U14328 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][6] ), .op(
        n12908) );
  nand2_1 U14329 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][6] ), .op(
        n12907) );
  nand2_1 U14330 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][6] ), .op(
        n12906) );
  nand2_1 U14331 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][6] ), .op(
        n12905) );
  nand2_1 U14332 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][6] ), .op(
        n12912) );
  nand2_1 U14333 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][6] ), .op(
        n12911) );
  nand2_1 U14334 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][6] ), .op(
        n12910) );
  nand2_1 U14335 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][6] ), .op(
        n12909) );
  nand2_1 U14336 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][6] ), .op(
        n12916) );
  nand2_1 U14337 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][6] ), .op(
        n12915) );
  nand2_1 U14338 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][6] ), .op(
        n12914) );
  nand2_1 U14339 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][6] ), .op(
        n12913) );
  nand2_1 U14340 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][6] ), .op(
        n12920) );
  nand2_1 U14341 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][6] ), .op(
        n12919) );
  nand2_1 U14342 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][6] ), .op(
        n12918) );
  nand2_1 U14343 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][6] ), .op(
        n12917) );
  mux2_1 U14344 ( .ip1(n18007), .ip2(n12929), .s(n14057), .op(n20485) );
  nand2_1 U14345 ( .ip1(n20485), .ip2(n13520), .op(n12931) );
  nand2_1 U14346 ( .ip1(n13521), .ip2(\pipeline/PC_DX [6]), .op(n12930) );
  nand2_1 U14347 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][6] ), .op(
        n12934) );
  nand2_1 U14348 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][6] ), .op(
        n12933) );
  nand2_1 U14349 ( .ip1(n12934), .ip2(n12933), .op(n12940) );
  nand2_1 U14350 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][6] ), .op(
        n12938) );
  nand2_1 U14351 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][6] ), .op(
        n12937) );
  nand2_1 U14352 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][6] ), .op(
        n12936) );
  nand2_1 U14353 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][6] ), .op(
        n12935) );
  not_ab_or_c_or_d U14354 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][6] ), 
        .ip3(n12940), .ip4(n12939), .op(n12972) );
  nand2_1 U14355 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][6] ), .op(
        n12944) );
  nand2_1 U14356 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][6] ), .op(
        n12943) );
  nand2_1 U14357 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][6] ), .op(
        n12942) );
  nand2_1 U14358 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][6] ), .op(
        n12941) );
  and4_1 U14359 ( .ip1(n12944), .ip2(n12943), .ip3(n12942), .ip4(n12941), .op(
        n12971) );
  nand2_1 U14360 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][6] ), .op(
        n12948) );
  nand2_1 U14361 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][6] ), .op(
        n12947) );
  nand2_1 U14362 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][6] ), .op(
        n12946) );
  nand2_1 U14363 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][6] ), .op(
        n12945) );
  and4_1 U14364 ( .ip1(n12948), .ip2(n12947), .ip3(n12946), .ip4(n12945), .op(
        n12970) );
  nand2_1 U14365 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][6] ), .op(
        n12952) );
  nand2_1 U14366 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][6] ), .op(
        n12951) );
  nand2_1 U14367 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][6] ), .op(
        n12950) );
  nand2_1 U14368 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][6] ), .op(
        n12949) );
  nand2_1 U14369 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][6] ), .op(
        n12956) );
  nand2_1 U14370 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][6] ), .op(
        n12955) );
  nand2_1 U14371 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][6] ), .op(
        n12954) );
  nand2_1 U14372 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][6] ), .op(
        n12953) );
  nand2_1 U14373 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][6] ), .op(
        n12960) );
  nand2_1 U14374 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][6] ), .op(
        n12959) );
  nand2_1 U14375 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][6] ), .op(
        n12958) );
  nand2_1 U14376 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][6] ), .op(
        n12957) );
  nand2_1 U14377 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][6] ), .op(
        n12964) );
  nand2_1 U14378 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][6] ), .op(
        n12963) );
  nand2_1 U14379 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][6] ), .op(
        n12962) );
  nand2_1 U14380 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][6] ), .op(
        n12961) );
  nand2_1 U14381 ( .ip1(n22065), .ip2(n10201), .op(n12975) );
  nand2_1 U14382 ( .ip1(n13445), .ip2(\pipeline/inst_DX [26]), .op(n12974) );
  nand2_1 U14383 ( .ip1(n12975), .ip2(n12974), .op(n17040) );
  nor2_1 U14384 ( .ip1(n17042), .ip2(n17040), .op(n13067) );
  nand2_1 U14385 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [7]), .op(n12978)
         );
  nand2_1 U14386 ( .ip1(\pipeline/alu_out_WB [7]), .ip2(n17895), .op(n12977)
         );
  nand2_1 U14387 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [7]), .op(
        n12976) );
  nand3_1 U14388 ( .ip1(n12978), .ip2(n12977), .ip3(n12976), .op(n18243) );
  nand2_1 U14389 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][7] ), .op(
        n12980) );
  nand2_1 U14390 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][7] ), .op(
        n12979) );
  nand2_1 U14391 ( .ip1(n12980), .ip2(n12979), .op(n12986) );
  nand2_1 U14392 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][7] ), .op(
        n12984) );
  nand2_1 U14393 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][7] ), .op(
        n12983) );
  nand2_1 U14394 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][7] ), .op(
        n12982) );
  nand2_1 U14395 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][7] ), .op(
        n12981) );
  not_ab_or_c_or_d U14396 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][7] ), 
        .ip3(n12986), .ip4(n12985), .op(n13018) );
  nand2_1 U14397 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][7] ), .op(
        n12990) );
  nand2_1 U14398 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][7] ), .op(
        n12989) );
  nand2_1 U14399 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][7] ), .op(
        n12988) );
  nand2_1 U14400 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][7] ), .op(
        n12987) );
  and4_1 U14401 ( .ip1(n12990), .ip2(n12989), .ip3(n12988), .ip4(n12987), .op(
        n13017) );
  nand2_1 U14402 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][7] ), .op(
        n12994) );
  nand2_1 U14403 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][7] ), .op(
        n12993) );
  nand2_1 U14404 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][7] ), .op(
        n12992) );
  nand2_1 U14405 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][7] ), .op(
        n12991) );
  and4_1 U14406 ( .ip1(n12994), .ip2(n12993), .ip3(n12992), .ip4(n12991), .op(
        n13016) );
  nand2_1 U14407 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][7] ), .op(
        n12998) );
  nand2_1 U14408 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][7] ), .op(
        n12997) );
  nand2_1 U14409 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][7] ), .op(
        n12996) );
  nand2_1 U14410 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][7] ), .op(
        n12995) );
  nand2_1 U14411 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][7] ), .op(
        n13002) );
  nand2_1 U14412 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][7] ), .op(
        n13001) );
  nand2_1 U14413 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][7] ), .op(
        n13000) );
  nand2_1 U14414 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][7] ), .op(
        n12999) );
  nand2_1 U14415 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][7] ), .op(
        n13006) );
  nand2_1 U14416 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][7] ), .op(
        n13005) );
  nand2_1 U14417 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][7] ), .op(
        n13004) );
  nand2_1 U14418 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][7] ), .op(
        n13003) );
  nand2_1 U14419 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][7] ), .op(
        n13010) );
  nand2_1 U14420 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][7] ), .op(
        n13009) );
  nand2_1 U14421 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][7] ), .op(
        n13008) );
  nand2_1 U14422 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][7] ), .op(
        n13007) );
  mux2_1 U14423 ( .ip1(n18243), .ip2(n13019), .s(n13162), .op(n15928) );
  nand2_1 U14424 ( .ip1(n15928), .ip2(n13520), .op(n13021) );
  nand2_1 U14425 ( .ip1(n13521), .ip2(\pipeline/PC_DX [7]), .op(n13020) );
  nand2_1 U14426 ( .ip1(n13445), .ip2(\pipeline/inst_DX [27]), .op(n13066) );
  nand2_1 U14427 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][7] ), .op(
        n13024) );
  nand2_1 U14428 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][7] ), .op(
        n13023) );
  nand2_1 U14429 ( .ip1(n13024), .ip2(n13023), .op(n13030) );
  nand2_1 U14430 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][7] ), .op(
        n13028) );
  nand2_1 U14431 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][7] ), .op(
        n13027) );
  nand2_1 U14432 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][7] ), .op(
        n13026) );
  nand2_1 U14433 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][7] ), .op(
        n13025) );
  not_ab_or_c_or_d U14434 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][7] ), 
        .ip3(n13030), .ip4(n13029), .op(n13062) );
  nand2_1 U14435 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][7] ), .op(
        n13034) );
  nand2_1 U14436 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][7] ), .op(
        n13033) );
  nand2_1 U14437 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][7] ), .op(
        n13032) );
  nand2_1 U14438 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][7] ), .op(
        n13031) );
  and4_1 U14439 ( .ip1(n13034), .ip2(n13033), .ip3(n13032), .ip4(n13031), .op(
        n13061) );
  nand2_1 U14440 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][7] ), .op(
        n13038) );
  nand2_1 U14441 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][7] ), .op(
        n13037) );
  nand2_1 U14442 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][7] ), .op(
        n13036) );
  nand2_1 U14443 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][7] ), .op(
        n13035) );
  and4_1 U14444 ( .ip1(n13038), .ip2(n13037), .ip3(n13036), .ip4(n13035), .op(
        n13060) );
  nand2_1 U14445 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][7] ), .op(
        n13042) );
  nand2_1 U14446 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][7] ), .op(
        n13041) );
  nand2_1 U14447 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][7] ), .op(
        n13040) );
  nand2_1 U14448 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][7] ), .op(
        n13039) );
  nand2_1 U14449 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][7] ), .op(
        n13046) );
  nand2_1 U14450 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][7] ), .op(
        n13045) );
  nand2_1 U14451 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][7] ), .op(
        n13044) );
  nand2_1 U14452 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][7] ), .op(
        n13043) );
  nand2_1 U14453 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][7] ), .op(
        n13050) );
  nand2_1 U14454 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][7] ), .op(
        n13049) );
  nand2_1 U14455 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][7] ), .op(
        n13048) );
  nand2_1 U14456 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][7] ), .op(
        n13047) );
  nand2_1 U14457 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][7] ), .op(
        n13054) );
  nand2_1 U14458 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][7] ), .op(
        n13053) );
  nand2_1 U14459 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][7] ), .op(
        n13052) );
  nand2_1 U14460 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][7] ), .op(
        n13051) );
  mux2_1 U14461 ( .ip1(n18243), .ip2(n13064), .s(n13063), .op(n17376) );
  nand2_1 U14462 ( .ip1(n17376), .ip2(n10201), .op(n13065) );
  nor2_1 U14463 ( .ip1(n13067), .ip2(n13538), .op(n13544) );
  nand2_1 U14464 ( .ip1(n13068), .ip2(n13544), .op(n13536) );
  nand2_1 U14465 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [3]), .op(n13071)
         );
  nand2_1 U14466 ( .ip1(\pipeline/alu_out_WB [3]), .ip2(n17895), .op(n13070)
         );
  nand2_1 U14467 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [3]), .op(
        n13069) );
  nand3_1 U14468 ( .ip1(n13071), .ip2(n13070), .ip3(n13069), .op(n17900) );
  nand2_1 U14469 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][3] ), .op(
        n13074) );
  nand2_1 U14470 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][3] ), .op(
        n13073) );
  nand2_1 U14471 ( .ip1(n13074), .ip2(n13073), .op(n13080) );
  nand2_1 U14472 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][3] ), .op(
        n13078) );
  nand2_1 U14473 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][3] ), .op(
        n13077) );
  nand2_1 U14474 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][3] ), .op(
        n13076) );
  nand2_1 U14475 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][3] ), .op(
        n13075) );
  not_ab_or_c_or_d U14476 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][3] ), 
        .ip3(n13080), .ip4(n13079), .op(n13112) );
  nand2_1 U14477 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][3] ), .op(
        n13084) );
  nand2_1 U14478 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][3] ), .op(
        n13083) );
  nand2_1 U14479 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][3] ), .op(
        n13082) );
  nand2_1 U14480 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][3] ), .op(
        n13081) );
  and4_1 U14481 ( .ip1(n13084), .ip2(n13083), .ip3(n13082), .ip4(n13081), .op(
        n13111) );
  nand2_1 U14482 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][3] ), .op(
        n13088) );
  nand2_1 U14483 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][3] ), .op(
        n13087) );
  nand2_1 U14484 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][3] ), .op(
        n13086) );
  nand2_1 U14485 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][3] ), .op(
        n13085) );
  and4_1 U14486 ( .ip1(n13088), .ip2(n13087), .ip3(n13086), .ip4(n13085), .op(
        n13110) );
  nand2_1 U14487 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][3] ), .op(
        n13092) );
  nand2_1 U14488 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][3] ), .op(
        n13091) );
  nand2_1 U14489 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][3] ), .op(
        n13090) );
  nand2_1 U14490 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][3] ), .op(
        n13089) );
  nand2_1 U14491 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][3] ), .op(
        n13096) );
  nand2_1 U14492 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][3] ), .op(
        n13095) );
  nand2_1 U14493 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][3] ), .op(
        n13094) );
  nand2_1 U14494 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][3] ), .op(
        n13093) );
  nand2_1 U14495 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][3] ), .op(
        n13100) );
  nand2_1 U14496 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][3] ), .op(
        n13099) );
  nand2_1 U14497 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][3] ), .op(
        n13098) );
  nand2_1 U14498 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][3] ), .op(
        n13097) );
  nand2_1 U14499 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][3] ), .op(
        n13104) );
  nand2_1 U14500 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][3] ), .op(
        n13103) );
  nand2_1 U14501 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][3] ), .op(
        n13102) );
  nand2_1 U14502 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][3] ), .op(
        n13101) );
  nand2_2 U14503 ( .ip1(n13115), .ip2(n13114), .op(n22059) );
  inv_1 U14504 ( .ip(\pipeline/inst_DX [10]), .op(n13116) );
  nor2_1 U14505 ( .ip1(n13443), .ip2(n13116), .op(n13119) );
  nor2_1 U14506 ( .ip1(n13117), .ip2(n13318), .op(n13118) );
  nor2_1 U14507 ( .ip1(n13119), .ip2(n13118), .op(n13120) );
  nand2_1 U14508 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][3] ), .op(
        n13123) );
  nand2_1 U14509 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][3] ), .op(
        n13122) );
  nand2_1 U14510 ( .ip1(n13123), .ip2(n13122), .op(n13129) );
  nand2_1 U14511 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][3] ), .op(
        n13127) );
  nand2_1 U14512 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][3] ), .op(
        n13126) );
  nand2_1 U14513 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][3] ), .op(
        n13125) );
  nand2_1 U14514 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][3] ), .op(
        n13124) );
  not_ab_or_c_or_d U14515 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][3] ), 
        .ip3(n13129), .ip4(n13128), .op(n13161) );
  nand2_1 U14516 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][3] ), .op(
        n13133) );
  nand2_1 U14517 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][3] ), .op(
        n13132) );
  nand2_1 U14518 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][3] ), .op(
        n13131) );
  nand2_1 U14519 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][3] ), .op(
        n13130) );
  and4_1 U14520 ( .ip1(n13133), .ip2(n13132), .ip3(n13131), .ip4(n13130), .op(
        n13160) );
  nand2_1 U14521 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][3] ), .op(
        n13137) );
  nand2_1 U14522 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][3] ), .op(
        n13136) );
  nand2_1 U14523 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][3] ), .op(
        n13135) );
  nand2_1 U14524 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][3] ), .op(
        n13134) );
  and4_1 U14525 ( .ip1(n13137), .ip2(n13136), .ip3(n13135), .ip4(n13134), .op(
        n13159) );
  nand2_1 U14526 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][3] ), .op(
        n13141) );
  nand2_1 U14527 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][3] ), .op(
        n13140) );
  nand2_1 U14528 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][3] ), .op(
        n13139) );
  nand2_1 U14529 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][3] ), .op(
        n13138) );
  nand2_1 U14530 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][3] ), .op(
        n13145) );
  nand2_1 U14531 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][3] ), .op(
        n13144) );
  nand2_1 U14532 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][3] ), .op(
        n13143) );
  nand2_1 U14533 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][3] ), .op(
        n13142) );
  nand2_1 U14534 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][3] ), .op(
        n13149) );
  nand2_1 U14535 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][3] ), .op(
        n13148) );
  nand2_1 U14536 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][3] ), .op(
        n13147) );
  nand2_1 U14537 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][3] ), .op(
        n13146) );
  nand2_1 U14538 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][3] ), .op(
        n13153) );
  nand2_1 U14539 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][3] ), .op(
        n13152) );
  nand2_1 U14540 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][3] ), .op(
        n13151) );
  nand2_1 U14541 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][3] ), .op(
        n13150) );
  mux2_1 U14542 ( .ip1(n17900), .ip2(n13163), .s(n13162), .op(n15796) );
  nand2_1 U14543 ( .ip1(n15796), .ip2(n13520), .op(n13165) );
  nand2_1 U14544 ( .ip1(n13521), .ip2(\pipeline/PC_DX [3]), .op(n13164) );
  nand2_1 U14545 ( .ip1(n16776), .ip2(n10195), .op(n13271) );
  nor2_1 U14546 ( .ip1(n16776), .ip2(n10195), .op(n13528) );
  nand2_1 U14547 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][2] ), .op(
        n13170) );
  nand2_1 U14548 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][2] ), .op(
        n13169) );
  nand2_1 U14549 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][2] ), .op(
        n13168) );
  nand2_1 U14550 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][2] ), .op(
        n13167) );
  and4_1 U14551 ( .ip1(n13170), .ip2(n13169), .ip3(n13168), .ip4(n13167), .op(
        n13174) );
  nand2_1 U14552 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][2] ), .op(
        n13173) );
  nand2_1 U14553 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][2] ), .op(
        n13172) );
  nand2_1 U14554 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][2] ), .op(
        n13171) );
  nand2_1 U14555 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][2] ), .op(
        n13178) );
  nand2_1 U14556 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][2] ), .op(
        n13177) );
  nand2_1 U14557 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][2] ), .op(
        n13176) );
  nand2_1 U14558 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][2] ), .op(
        n13175) );
  nand2_1 U14559 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][2] ), .op(
        n13182) );
  nand2_1 U14560 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][2] ), .op(
        n13181) );
  nand2_1 U14561 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][2] ), .op(
        n13180) );
  nand2_1 U14562 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][2] ), .op(
        n13179) );
  nand2_1 U14563 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][2] ), .op(
        n13186) );
  nand2_1 U14564 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][2] ), .op(
        n13185) );
  nand2_1 U14565 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][2] ), .op(
        n13184) );
  nand2_1 U14566 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][2] ), .op(
        n13183) );
  nand2_1 U14567 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][2] ), .op(
        n13190) );
  nand2_1 U14568 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][2] ), .op(
        n13189) );
  nand2_1 U14569 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][2] ), .op(
        n13188) );
  nand2_1 U14570 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][2] ), .op(
        n13187) );
  nand2_1 U14571 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][2] ), .op(
        n13194) );
  nand2_1 U14572 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][2] ), .op(
        n13193) );
  nand2_1 U14573 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][2] ), .op(
        n13192) );
  nand2_1 U14574 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][2] ), .op(
        n13191) );
  nand2_1 U14575 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][2] ), .op(
        n13198) );
  nand2_1 U14576 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][2] ), .op(
        n13197) );
  nand2_1 U14577 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][2] ), .op(
        n13196) );
  nand2_1 U14578 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][2] ), .op(
        n13195) );
  or4_1 U14579 ( .ip1(n13202), .ip2(n13201), .ip3(n13200), .ip4(n13199), .op(
        n13203) );
  nor2_1 U14580 ( .ip1(n15290), .ip2(n13220), .op(n13215) );
  nor2_1 U14581 ( .ip1(n13207), .ip2(n13318), .op(n13214) );
  inv_1 U14582 ( .ip(n13443), .op(n13208) );
  nand2_1 U14583 ( .ip1(n13208), .ip2(\pipeline/inst_DX [9]), .op(n13212) );
  nand2_1 U14584 ( .ip1(n13210), .ip2(n13209), .op(n13211) );
  nand2_1 U14585 ( .ip1(n13212), .ip2(n13211), .op(n13213) );
  not_ab_or_c_or_d U14586 ( .ip1(n13315), .ip2(n13215), .ip3(n13214), .ip4(
        n13213), .op(n13223) );
  inv_1 U14587 ( .ip(\pipeline/alu_out_WB [2]), .op(n13216) );
  nor2_1 U14588 ( .ip1(\pipeline/wb_src_sel_WB [1]), .ip2(n13216), .op(n13219)
         );
  inv_1 U14589 ( .ip(\pipeline/md_resp_result [2]), .op(n14920) );
  nor2_1 U14590 ( .ip1(n13217), .ip2(n14920), .op(n13218) );
  not_ab_or_c_or_d U14591 ( .ip1(\pipeline/csr_rdata_WB [2]), .ip2(n13368), 
        .ip3(n13219), .ip4(n13218), .op(n15291) );
  nor2_1 U14592 ( .ip1(n15291), .ip2(n13220), .op(n13221) );
  nand2_1 U14593 ( .ip1(n12880), .ip2(n13221), .op(n13222) );
  nand2_1 U14594 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][2] ), .op(
        n13225) );
  nand2_1 U14595 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][2] ), .op(
        n13224) );
  nand2_1 U14596 ( .ip1(n13225), .ip2(n13224), .op(n13231) );
  nand2_1 U14597 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][2] ), .op(
        n13229) );
  nand2_1 U14598 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][2] ), .op(
        n13228) );
  nand2_1 U14599 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][2] ), .op(
        n13227) );
  nand2_1 U14600 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][2] ), .op(
        n13226) );
  not_ab_or_c_or_d U14601 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][2] ), 
        .ip3(n13231), .ip4(n13230), .op(n13263) );
  nand2_1 U14602 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][2] ), .op(
        n13235) );
  nand2_1 U14603 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][2] ), .op(
        n13234) );
  nand2_1 U14604 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][2] ), .op(
        n13233) );
  nand2_1 U14605 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][2] ), .op(
        n13232) );
  and4_1 U14606 ( .ip1(n13235), .ip2(n13234), .ip3(n13233), .ip4(n13232), .op(
        n13262) );
  nand2_1 U14607 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][2] ), .op(
        n13239) );
  nand2_1 U14608 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][2] ), .op(
        n13238) );
  nand2_1 U14609 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][2] ), .op(
        n13237) );
  nand2_1 U14610 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][2] ), .op(
        n13236) );
  and4_1 U14611 ( .ip1(n13239), .ip2(n13238), .ip3(n13237), .ip4(n13236), .op(
        n13261) );
  nand2_1 U14612 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][2] ), .op(
        n13243) );
  nand2_1 U14613 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][2] ), .op(
        n13242) );
  nand2_1 U14614 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][2] ), .op(
        n13241) );
  nand2_1 U14615 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][2] ), .op(
        n13240) );
  nand2_1 U14616 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][2] ), .op(
        n13247) );
  nand2_1 U14617 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][2] ), .op(
        n13246) );
  nand2_1 U14618 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][2] ), .op(
        n13245) );
  nand2_1 U14619 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][2] ), .op(
        n13244) );
  nand2_1 U14620 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][2] ), .op(
        n13251) );
  nand2_1 U14621 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][2] ), .op(
        n13250) );
  nand2_1 U14622 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][2] ), .op(
        n13249) );
  nand2_1 U14623 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][2] ), .op(
        n13248) );
  nand2_1 U14624 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][2] ), .op(
        n13255) );
  nand2_1 U14625 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][2] ), .op(
        n13254) );
  nand2_1 U14626 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][2] ), .op(
        n13253) );
  nand2_1 U14627 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][2] ), .op(
        n13252) );
  inv_1 U14628 ( .ip(n15291), .op(n21155) );
  nand2_1 U14629 ( .ip1(n13521), .ip2(\pipeline/PC_DX [2]), .op(n13267) );
  nand2_1 U14630 ( .ip1(n10198), .ip2(n13728), .op(n13269) );
  or2_1 U14631 ( .ip1(n13528), .ip2(n13269), .op(n13270) );
  nand2_1 U14632 ( .ip1(n13271), .ip2(n13270), .op(n13534) );
  nand2_1 U14633 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [1]), .op(n13274)
         );
  nand2_1 U14634 ( .ip1(\pipeline/alu_out_WB [1]), .ip2(n17895), .op(n13273)
         );
  nand2_1 U14635 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [1]), .op(
        n13272) );
  nand3_1 U14636 ( .ip1(n13274), .ip2(n13273), .ip3(n13272), .op(n18016) );
  nand2_1 U14637 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][1] ), .op(
        n13276) );
  nand2_1 U14638 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][1] ), .op(
        n13275) );
  nand2_1 U14639 ( .ip1(n13276), .ip2(n13275), .op(n13282) );
  nand2_1 U14640 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][1] ), .op(
        n13280) );
  nand2_1 U14641 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][1] ), .op(
        n13279) );
  nand2_1 U14642 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][1] ), .op(
        n13278) );
  nand2_1 U14643 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][1] ), .op(
        n13277) );
  not_ab_or_c_or_d U14644 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][1] ), 
        .ip3(n13282), .ip4(n13281), .op(n13314) );
  nand2_1 U14645 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][1] ), .op(
        n13286) );
  nand2_1 U14646 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][1] ), .op(
        n13285) );
  nand2_1 U14647 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][1] ), .op(
        n13284) );
  nand2_1 U14648 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][1] ), .op(
        n13283) );
  and4_1 U14649 ( .ip1(n13286), .ip2(n13285), .ip3(n13284), .ip4(n13283), .op(
        n13313) );
  nand2_1 U14650 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][1] ), .op(
        n13290) );
  nand2_1 U14651 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][1] ), .op(
        n13289) );
  nand2_1 U14652 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][1] ), .op(
        n13288) );
  nand2_1 U14653 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][1] ), .op(
        n13287) );
  and4_1 U14654 ( .ip1(n13290), .ip2(n13289), .ip3(n13288), .ip4(n13287), .op(
        n13312) );
  nand2_1 U14655 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][1] ), .op(
        n13294) );
  nand2_1 U14656 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][1] ), .op(
        n13293) );
  nand2_1 U14657 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][1] ), .op(
        n13292) );
  nand2_1 U14658 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][1] ), .op(
        n13291) );
  nand2_1 U14659 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][1] ), .op(
        n13298) );
  nand2_1 U14660 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][1] ), .op(
        n13297) );
  nand2_1 U14661 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][1] ), .op(
        n13296) );
  nand2_1 U14662 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][1] ), .op(
        n13295) );
  nand2_1 U14663 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][1] ), .op(
        n13302) );
  nand2_1 U14664 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][1] ), .op(
        n13301) );
  nand2_1 U14665 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][1] ), .op(
        n13300) );
  nand2_1 U14666 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][1] ), .op(
        n13299) );
  nand2_1 U14667 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][1] ), .op(
        n13306) );
  nand2_1 U14668 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][1] ), .op(
        n13305) );
  nand2_1 U14669 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][1] ), .op(
        n13304) );
  nand2_1 U14670 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][1] ), .op(
        n13303) );
  mux2_1 U14671 ( .ip1(n18016), .ip2(n13316), .s(n13315), .op(n22055) );
  nand2_1 U14672 ( .ip1(n22055), .ip2(n10201), .op(n13323) );
  inv_1 U14673 ( .ip(\pipeline/inst_DX [8]), .op(n13317) );
  nor2_1 U14674 ( .ip1(n13443), .ip2(n13317), .op(n13321) );
  nor2_1 U14675 ( .ip1(n13319), .ip2(n13318), .op(n13320) );
  nor2_1 U14676 ( .ip1(n13321), .ip2(n13320), .op(n13322) );
  nand2_1 U14677 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][1] ), .op(
        n13325) );
  nand2_1 U14678 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][1] ), .op(
        n13324) );
  nand2_1 U14679 ( .ip1(n13325), .ip2(n13324), .op(n13331) );
  nand2_1 U14680 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][1] ), .op(
        n13329) );
  nand2_1 U14681 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][1] ), .op(
        n13328) );
  nand2_1 U14682 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][1] ), .op(
        n13327) );
  nand2_1 U14683 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][1] ), .op(
        n13326) );
  not_ab_or_c_or_d U14684 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][1] ), 
        .ip3(n13331), .ip4(n13330), .op(n13363) );
  nand2_1 U14685 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][1] ), .op(
        n13335) );
  nand2_1 U14686 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][1] ), .op(
        n13334) );
  nand2_1 U14687 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][1] ), .op(
        n13333) );
  nand2_1 U14688 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][1] ), .op(
        n13332) );
  and4_1 U14689 ( .ip1(n13335), .ip2(n13334), .ip3(n13333), .ip4(n13332), .op(
        n13362) );
  nand2_1 U14690 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][1] ), .op(
        n13339) );
  nand2_1 U14691 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][1] ), .op(
        n13338) );
  nand2_1 U14692 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][1] ), .op(
        n13337) );
  nand2_1 U14693 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][1] ), .op(
        n13336) );
  and4_1 U14694 ( .ip1(n13339), .ip2(n13338), .ip3(n13337), .ip4(n13336), .op(
        n13361) );
  nand2_1 U14695 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][1] ), .op(
        n13343) );
  nand2_1 U14696 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][1] ), .op(
        n13342) );
  nand2_1 U14697 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][1] ), .op(
        n13341) );
  nand2_1 U14698 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][1] ), .op(
        n13340) );
  nand2_1 U14699 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][1] ), .op(
        n13347) );
  nand2_1 U14700 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][1] ), .op(
        n13346) );
  nand2_1 U14701 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][1] ), .op(
        n13345) );
  nand2_1 U14702 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][1] ), .op(
        n13344) );
  nand2_1 U14703 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][1] ), .op(
        n13351) );
  nand2_1 U14704 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][1] ), .op(
        n13350) );
  nand2_1 U14705 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][1] ), .op(
        n13349) );
  nand2_1 U14706 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][1] ), .op(
        n13348) );
  nand2_1 U14707 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][1] ), .op(
        n13355) );
  nand2_1 U14708 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][1] ), .op(
        n13354) );
  nand2_1 U14709 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][1] ), .op(
        n13353) );
  nand2_1 U14710 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][1] ), .op(
        n13352) );
  mux2_1 U14711 ( .ip1(n18016), .ip2(n13365), .s(n13364), .op(n14597) );
  nand2_1 U14712 ( .ip1(n14597), .ip2(n13520), .op(n13367) );
  nand2_1 U14713 ( .ip1(n13521), .ip2(\pipeline/PC_DX [1]), .op(n13366) );
  nand2_1 U14714 ( .ip1(n13525), .ip2(n16608), .op(n13722) );
  nand2_1 U14715 ( .ip1(n13368), .ip2(\pipeline/csr_rdata_WB [0]), .op(n13372)
         );
  nand2_1 U14716 ( .ip1(\pipeline/alu_out_WB [0]), .ip2(n17895), .op(n13371)
         );
  nand2_1 U14717 ( .ip1(n13369), .ip2(\pipeline/md_resp_result [0]), .op(
        n13370) );
  nand3_1 U14718 ( .ip1(n13372), .ip2(n13371), .ip3(n13370), .op(n21239) );
  nand2_1 U14719 ( .ip1(n22097), .ip2(\pipeline/regfile/data[4][0] ), .op(
        n13374) );
  nand2_1 U14720 ( .ip1(n22109), .ip2(\pipeline/regfile/data[1][0] ), .op(
        n13373) );
  nand2_1 U14721 ( .ip1(n13374), .ip2(n13373), .op(n13383) );
  nand2_1 U14722 ( .ip1(n15338), .ip2(\pipeline/regfile/data[2][0] ), .op(
        n13381) );
  nand2_1 U14723 ( .ip1(n13375), .ip2(\pipeline/regfile/data[16][0] ), .op(
        n13380) );
  nand2_1 U14724 ( .ip1(n13376), .ip2(\pipeline/regfile/data[3][0] ), .op(
        n13379) );
  nand2_1 U14725 ( .ip1(n13377), .ip2(\pipeline/regfile/data[20][0] ), .op(
        n13378) );
  not_ab_or_c_or_d U14726 ( .ip1(n13384), .ip2(\pipeline/regfile/data[14][0] ), 
        .ip3(n13383), .ip4(n13382), .op(n13440) );
  nand2_1 U14727 ( .ip1(n13385), .ip2(\pipeline/regfile/data[9][0] ), .op(
        n13392) );
  nand2_1 U14728 ( .ip1(n13386), .ip2(\pipeline/regfile/data[21][0] ), .op(
        n13391) );
  nand2_1 U14729 ( .ip1(n13387), .ip2(\pipeline/regfile/data[24][0] ), .op(
        n13390) );
  nand2_1 U14730 ( .ip1(n13388), .ip2(\pipeline/regfile/data[10][0] ), .op(
        n13389) );
  and4_1 U14731 ( .ip1(n13392), .ip2(n13391), .ip3(n13390), .ip4(n13389), .op(
        n13439) );
  nand2_1 U14732 ( .ip1(n13393), .ip2(\pipeline/regfile/data[7][0] ), .op(
        n13400) );
  nand2_1 U14733 ( .ip1(n13394), .ip2(\pipeline/regfile/data[8][0] ), .op(
        n13399) );
  nand2_1 U14734 ( .ip1(n13395), .ip2(\pipeline/regfile/data[23][0] ), .op(
        n13398) );
  nand2_1 U14735 ( .ip1(n13396), .ip2(\pipeline/regfile/data[17][0] ), .op(
        n13397) );
  and4_1 U14736 ( .ip1(n13400), .ip2(n13399), .ip3(n13398), .ip4(n13397), .op(
        n13438) );
  nand2_1 U14737 ( .ip1(n13401), .ip2(\pipeline/regfile/data[11][0] ), .op(
        n13408) );
  nand2_1 U14738 ( .ip1(n13402), .ip2(\pipeline/regfile/data[25][0] ), .op(
        n13407) );
  nand2_1 U14739 ( .ip1(n13403), .ip2(\pipeline/regfile/data[18][0] ), .op(
        n13406) );
  nand2_1 U14740 ( .ip1(n13404), .ip2(\pipeline/regfile/data[19][0] ), .op(
        n13405) );
  nand2_1 U14741 ( .ip1(n13409), .ip2(\pipeline/regfile/data[6][0] ), .op(
        n13416) );
  nand2_1 U14742 ( .ip1(n13410), .ip2(\pipeline/regfile/data[27][0] ), .op(
        n13415) );
  nand2_1 U14743 ( .ip1(n13411), .ip2(\pipeline/regfile/data[26][0] ), .op(
        n13414) );
  nand2_1 U14744 ( .ip1(n13412), .ip2(\pipeline/regfile/data[22][0] ), .op(
        n13413) );
  nand2_1 U14745 ( .ip1(n13417), .ip2(\pipeline/regfile/data[15][0] ), .op(
        n13424) );
  nand2_1 U14746 ( .ip1(n13418), .ip2(\pipeline/regfile/data[5][0] ), .op(
        n13423) );
  nand2_1 U14747 ( .ip1(n13419), .ip2(\pipeline/regfile/data[12][0] ), .op(
        n13422) );
  nand2_1 U14748 ( .ip1(n13420), .ip2(\pipeline/regfile/data[13][0] ), .op(
        n13421) );
  nand2_1 U14749 ( .ip1(n13425), .ip2(\pipeline/regfile/data[30][0] ), .op(
        n13432) );
  nand2_1 U14750 ( .ip1(n13426), .ip2(\pipeline/regfile/data[28][0] ), .op(
        n13431) );
  nand2_1 U14751 ( .ip1(n13427), .ip2(\pipeline/regfile/data[31][0] ), .op(
        n13430) );
  nand2_1 U14752 ( .ip1(n13428), .ip2(\pipeline/regfile/data[29][0] ), .op(
        n13429) );
  mux2_1 U14753 ( .ip1(n21239), .ip2(n13442), .s(n13441), .op(n22053) );
  nand2_1 U14754 ( .ip1(n22053), .ip2(n10201), .op(n13447) );
  mux2_1 U14755 ( .ip1(\pipeline/inst_DX [7]), .ip2(\pipeline/inst_DX [20]), 
        .s(n13443), .op(n13444) );
  nand2_1 U14756 ( .ip1(n13445), .ip2(n13444), .op(n13446) );
  nand2_1 U14757 ( .ip1(n13447), .ip2(n13446), .op(n16487) );
  nand2_1 U14758 ( .ip1(n13448), .ip2(\pipeline/regfile/data[8][0] ), .op(
        n13451) );
  nand2_1 U14759 ( .ip1(n13449), .ip2(\pipeline/regfile/data[10][0] ), .op(
        n13450) );
  nand2_1 U14760 ( .ip1(n13451), .ip2(n13450), .op(n13461) );
  nand2_1 U14761 ( .ip1(n13452), .ip2(\pipeline/regfile/data[21][0] ), .op(
        n13459) );
  nand2_1 U14762 ( .ip1(n13453), .ip2(\pipeline/regfile/data[17][0] ), .op(
        n13458) );
  nand2_1 U14763 ( .ip1(n13454), .ip2(\pipeline/regfile/data[7][0] ), .op(
        n13457) );
  nand2_1 U14764 ( .ip1(n13455), .ip2(\pipeline/regfile/data[1][0] ), .op(
        n13456) );
  not_ab_or_c_or_d U14765 ( .ip1(n13462), .ip2(\pipeline/regfile/data[28][0] ), 
        .ip3(n13461), .ip4(n13460), .op(n13518) );
  nand2_1 U14766 ( .ip1(n13463), .ip2(\pipeline/regfile/data[27][0] ), .op(
        n13470) );
  nand2_1 U14767 ( .ip1(n13464), .ip2(\pipeline/regfile/data[9][0] ), .op(
        n13469) );
  nand2_1 U14768 ( .ip1(n13465), .ip2(\pipeline/regfile/data[2][0] ), .op(
        n13468) );
  nand2_1 U14769 ( .ip1(n13466), .ip2(\pipeline/regfile/data[26][0] ), .op(
        n13467) );
  and4_1 U14770 ( .ip1(n13470), .ip2(n13469), .ip3(n13468), .ip4(n13467), .op(
        n13517) );
  nand2_1 U14771 ( .ip1(n13471), .ip2(\pipeline/regfile/data[16][0] ), .op(
        n13478) );
  nand2_1 U14772 ( .ip1(n13472), .ip2(\pipeline/regfile/data[4][0] ), .op(
        n13477) );
  nand2_1 U14773 ( .ip1(n13473), .ip2(\pipeline/regfile/data[24][0] ), .op(
        n13476) );
  nand2_1 U14774 ( .ip1(n13474), .ip2(\pipeline/regfile/data[20][0] ), .op(
        n13475) );
  and4_1 U14775 ( .ip1(n13478), .ip2(n13477), .ip3(n13476), .ip4(n13475), .op(
        n13516) );
  nand2_1 U14776 ( .ip1(n13479), .ip2(\pipeline/regfile/data[25][0] ), .op(
        n13486) );
  nand2_1 U14777 ( .ip1(n13480), .ip2(\pipeline/regfile/data[3][0] ), .op(
        n13485) );
  nand2_1 U14778 ( .ip1(n13481), .ip2(\pipeline/regfile/data[6][0] ), .op(
        n13484) );
  nand2_1 U14779 ( .ip1(n13482), .ip2(\pipeline/regfile/data[5][0] ), .op(
        n13483) );
  nand2_1 U14780 ( .ip1(n13487), .ip2(\pipeline/regfile/data[18][0] ), .op(
        n13494) );
  nand2_1 U14781 ( .ip1(n13488), .ip2(\pipeline/regfile/data[23][0] ), .op(
        n13493) );
  nand2_1 U14782 ( .ip1(n13489), .ip2(\pipeline/regfile/data[11][0] ), .op(
        n13492) );
  nand2_1 U14783 ( .ip1(n13490), .ip2(\pipeline/regfile/data[19][0] ), .op(
        n13491) );
  nand2_1 U14784 ( .ip1(n13495), .ip2(\pipeline/regfile/data[29][0] ), .op(
        n13502) );
  nand2_1 U14785 ( .ip1(n13496), .ip2(\pipeline/regfile/data[22][0] ), .op(
        n13501) );
  nand2_1 U14786 ( .ip1(n13497), .ip2(\pipeline/regfile/data[15][0] ), .op(
        n13500) );
  nand2_1 U14787 ( .ip1(n13498), .ip2(\pipeline/regfile/data[31][0] ), .op(
        n13499) );
  nand2_1 U14788 ( .ip1(n13503), .ip2(\pipeline/regfile/data[14][0] ), .op(
        n13510) );
  nand2_1 U14789 ( .ip1(n13504), .ip2(\pipeline/regfile/data[13][0] ), .op(
        n13509) );
  nand2_1 U14790 ( .ip1(n13505), .ip2(\pipeline/regfile/data[30][0] ), .op(
        n13508) );
  nand2_1 U14791 ( .ip1(n13506), .ip2(\pipeline/regfile/data[12][0] ), .op(
        n13507) );
  mux2_1 U14792 ( .ip1(n21239), .ip2(n13519), .s(n13162), .op(n18022) );
  nand2_1 U14793 ( .ip1(n18022), .ip2(n13520), .op(n13523) );
  nand2_1 U14794 ( .ip1(n13521), .ip2(\pipeline/PC_DX [0]), .op(n13522) );
  nand2_1 U14795 ( .ip1(n16487), .ip2(n13870), .op(n13804) );
  inv_1 U14796 ( .ip(n13807), .op(n16732) );
  nor2_1 U14797 ( .ip1(n16732), .ip2(n16608), .op(n13526) );
  or2_1 U14798 ( .ip1(n13804), .ip2(n13526), .op(n13527) );
  nand2_1 U14799 ( .ip1(n13722), .ip2(n13527), .op(n13531) );
  nor2_1 U14800 ( .ip1(n10198), .ip2(n13728), .op(n13529) );
  nor2_1 U14801 ( .ip1(n13529), .ip2(n13528), .op(n13530) );
  nand2_1 U14802 ( .ip1(n13531), .ip2(n13530), .op(n13532) );
  inv_1 U14803 ( .ip(n13532), .op(n13533) );
  nor2_1 U14804 ( .ip1(n13534), .ip2(n13533), .op(n13535) );
  or2_1 U14805 ( .ip1(n13536), .ip2(n13535), .op(n13549) );
  or2_1 U14806 ( .ip1(n13930), .ip2(n13538), .op(n13539) );
  nand2_1 U14807 ( .ip1(n13932), .ip2(n13539), .op(n13547) );
  nand2_1 U14808 ( .ip1(n13540), .ip2(n17199), .op(n13542) );
  or2_1 U14809 ( .ip1(n13542), .ip2(n13541), .op(n13543) );
  nand2_1 U14810 ( .ip1(n13933), .ip2(n13543), .op(n13545) );
  and2_1 U14811 ( .ip1(n13545), .ip2(n13544), .op(n13546) );
  nor2_1 U14812 ( .ip1(n13547), .ip2(n13546), .op(n13548) );
  nand2_1 U14813 ( .ip1(n13549), .ip2(n13548), .op(n13550) );
  nand2_1 U14814 ( .ip1(n13551), .ip2(n13550), .op(n13565) );
  nand2_1 U14815 ( .ip1(n13552), .ip2(n16690), .op(n13556) );
  nand2_1 U14816 ( .ip1(n13553), .ip2(n16972), .op(n13924) );
  or2_1 U14817 ( .ip1(n13924), .ip2(n13554), .op(n13555) );
  nand2_1 U14818 ( .ip1(n13556), .ip2(n13555), .op(n13562) );
  inv_1 U14819 ( .ip(n13922), .op(n13557) );
  nand2_1 U14820 ( .ip1(n13557), .ip2(n13860), .op(n13558) );
  nand2_1 U14821 ( .ip1(n10206), .ip2(n17457), .op(n13921) );
  nand2_1 U14822 ( .ip1(n13558), .ip2(n13921), .op(n13560) );
  and2_1 U14823 ( .ip1(n13560), .ip2(n13559), .op(n13561) );
  nor2_1 U14824 ( .ip1(n13562), .ip2(n13561), .op(n13563) );
  or2_1 U14825 ( .ip1(n13563), .ip2(n13832), .op(n13564) );
  nand3_1 U14826 ( .ip1(n13833), .ip2(n13565), .ip3(n13564), .op(n13573) );
  nor2_1 U14827 ( .ip1(n13868), .ip2(n16418), .op(n13961) );
  inv_1 U14828 ( .ip(n13885), .op(n13955) );
  nor2_1 U14829 ( .ip1(n13961), .ip2(n13955), .op(n13567) );
  nand2_1 U14830 ( .ip1(n13567), .ip2(n13566), .op(n13568) );
  nor2_1 U14831 ( .ip1(n13569), .ip2(n13568), .op(n13571) );
  nand2_1 U14832 ( .ip1(n13573), .ip2(n13572), .op(n13574) );
  nand4_1 U14833 ( .ip1(n17786), .ip2(dmem_hsize[0]), .ip3(n13577), .ip4(
        n13576), .op(n13754) );
  inv_1 U14834 ( .ip(n16477), .op(n13580) );
  nand2_1 U14835 ( .ip1(n17786), .ip2(n13580), .op(n13592) );
  inv_1 U14836 ( .ip(n13592), .op(n13589) );
  nand2_1 U14837 ( .ip1(n15312), .ip2(n17765), .op(n13581) );
  nand2_1 U14838 ( .ip1(dmem_hsize[1]), .ip2(n13581), .op(n13587) );
  nand2_1 U14839 ( .ip1(n14596), .ip2(n13582), .op(n13584) );
  nand2_1 U14840 ( .ip1(dmem_hsize[0]), .ip2(\pipeline/dmem_type[2] ), .op(
        n13583) );
  nand2_1 U14841 ( .ip1(n13584), .ip2(n13583), .op(n13585) );
  nand2_1 U14842 ( .ip1(\pipeline/inst_DX [30]), .ip2(n13585), .op(n13586) );
  nand2_1 U14843 ( .ip1(n13587), .ip2(n13586), .op(n13588) );
  nand2_1 U14844 ( .ip1(n13589), .ip2(n13588), .op(n13591) );
  nor3_1 U14845 ( .ip1(n16479), .ip2(n16483), .ip3(n17765), .op(n13595) );
  nand2_1 U14846 ( .ip1(dmem_hsize[1]), .ip2(n13595), .op(n13590) );
  nand2_1 U14847 ( .ip1(n13591), .ip2(n13590), .op(n16913) );
  nor3_1 U14848 ( .ip1(dmem_hsize[1]), .ip2(n15308), .ip3(n15312), .op(n13593)
         );
  nor3_1 U14849 ( .ip1(n16478), .ip2(n13593), .ip3(n13592), .op(n13594) );
  nor2_1 U14850 ( .ip1(n13595), .ip2(n13594), .op(n13895) );
  nor2_1 U14851 ( .ip1(n13895), .ip2(n13754), .op(n16525) );
  inv_1 U14852 ( .ip(n13596), .op(n20856) );
  nand2_1 U14853 ( .ip1(n20856), .ip2(n10196), .op(n13610) );
  or2_1 U14854 ( .ip1(n20856), .ip2(n10196), .op(n13746) );
  inv_1 U14855 ( .ip(n11935), .op(n13597) );
  nand2_1 U14856 ( .ip1(n13600), .ip2(n13599), .op(n13975) );
  inv_1 U14857 ( .ip(n13742), .op(n16533) );
  or2_1 U14858 ( .ip1(n16533), .ip2(n13601), .op(n13985) );
  nand2_1 U14859 ( .ip1(n11945), .ip2(n13779), .op(n13602) );
  inv_1 U14860 ( .ip(n10180), .op(n19068) );
  nand2_1 U14861 ( .ip1(n19067), .ip2(n19068), .op(n13984) );
  nand2_1 U14862 ( .ip1(n13602), .ip2(n13984), .op(n13603) );
  nand2_1 U14863 ( .ip1(n13977), .ip2(n13603), .op(n13604) );
  nand2_1 U14864 ( .ip1(n13975), .ip2(n13604), .op(n13605) );
  inv_1 U14865 ( .ip(n16550), .op(n17277) );
  nor2_1 U14866 ( .ip1(n17277), .ip2(n13665), .op(n13667) );
  inv_1 U14867 ( .ip(n13667), .op(n13616) );
  inv_1 U14868 ( .ip(n13614), .op(n13615) );
  nand2_1 U14869 ( .ip1(n16545), .ip2(n10192), .op(n13758) );
  nand2_1 U14870 ( .ip1(n13615), .ip2(n13758), .op(n14001) );
  nor2_1 U14871 ( .ip1(n10197), .ip2(n10188), .op(n13908) );
  nand2_1 U14872 ( .ip1(n16935), .ip2(n10178), .op(n13845) );
  nand2_1 U14873 ( .ip1(n16594), .ip2(n13654), .op(n13884) );
  inv_1 U14874 ( .ip(n18731), .op(n18730) );
  nor2_1 U14875 ( .ip1(n18730), .ip2(n10186), .op(n13655) );
  inv_1 U14876 ( .ip(n13655), .op(n13620) );
  nand2_1 U14877 ( .ip1(n13884), .ip2(n13620), .op(n13621) );
  inv_1 U14878 ( .ip(n13947), .op(n13886) );
  nand2_1 U14879 ( .ip1(n13886), .ip2(n13954), .op(n13642) );
  inv_1 U14880 ( .ip(n13948), .op(n13624) );
  or2_1 U14881 ( .ip1(n19430), .ip2(n16846), .op(n13623) );
  nand2_1 U14882 ( .ip1(n13624), .ip2(n13623), .op(n13625) );
  nor2_1 U14883 ( .ip1(n13642), .ip2(n13625), .op(n13685) );
  inv_1 U14884 ( .ip(n20728), .op(n20727) );
  nand2_1 U14885 ( .ip1(n20727), .ip2(n16838), .op(n13628) );
  inv_1 U14886 ( .ip(n17142), .op(n17143) );
  nand2_1 U14887 ( .ip1(n17143), .ip2(n12138), .op(n13631) );
  inv_1 U14888 ( .ip(n13631), .op(n13633) );
  inv_1 U14889 ( .ip(n13636), .op(n19433) );
  inv_1 U14890 ( .ip(n13868), .op(n16845) );
  nand2_1 U14891 ( .ip1(n16498), .ip2(n16845), .op(n13638) );
  inv_1 U14892 ( .ip(n13638), .op(n13639) );
  nor2_1 U14893 ( .ip1(n13640), .ip2(n13639), .op(n13641) );
  nor2_1 U14894 ( .ip1(n13642), .ip2(n13641), .op(n13648) );
  inv_1 U14895 ( .ip(n16557), .op(n16855) );
  nand2_1 U14896 ( .ip1(n16855), .ip2(n16854), .op(n13956) );
  inv_1 U14897 ( .ip(n13956), .op(n13646) );
  or2_1 U14898 ( .ip1(n16559), .ip2(n16526), .op(n13644) );
  nor2_1 U14899 ( .ip1(n13644), .ip2(n13643), .op(n13645) );
  or2_1 U14900 ( .ip1(n13646), .ip2(n13645), .op(n13647) );
  not_ab_or_c_or_d U14901 ( .ip1(n13685), .ip2(n13959), .ip3(n13648), .ip4(
        n13647), .op(n13649) );
  or2_1 U14902 ( .ip1(n13686), .ip2(n13649), .op(n13741) );
  inv_1 U14903 ( .ip(n16935), .op(n16933) );
  inv_1 U14904 ( .ip(n10178), .op(n19051) );
  inv_1 U14905 ( .ip(n13845), .op(n13902) );
  nor2_1 U14906 ( .ip1(n13994), .ip2(n13902), .op(n13652) );
  nor2_1 U14907 ( .ip1(n13650), .ip2(n13652), .op(n13661) );
  inv_1 U14908 ( .ip(n13653), .op(n13659) );
  nor2_1 U14909 ( .ip1(n13993), .ip2(n13655), .op(n13657) );
  nand2_1 U14910 ( .ip1(n18730), .ip2(n10186), .op(n13992) );
  inv_1 U14911 ( .ip(n13992), .op(n13765) );
  inv_1 U14912 ( .ip(n17173), .op(n17171) );
  nand2_1 U14913 ( .ip1(n17171), .ip2(n18737), .op(n13854) );
  inv_1 U14914 ( .ip(n13854), .op(n13664) );
  inv_1 U14915 ( .ip(n16545), .op(n17531) );
  nand2_1 U14916 ( .ip1(n13662), .ip2(n17531), .op(n13855) );
  nor2_1 U14917 ( .ip1(n13614), .ip2(n13855), .op(n13663) );
  nor2_1 U14918 ( .ip1(n13664), .ip2(n13663), .op(n14005) );
  nand2_1 U14919 ( .ip1(n17277), .ip2(n13665), .op(n13996) );
  inv_1 U14920 ( .ip(n13996), .op(n13669) );
  nand2_1 U14921 ( .ip1(n14002), .ip2(n10236), .op(n13670) );
  nand2_1 U14922 ( .ip1(n14005), .ip2(n13670), .op(n13672) );
  nand2_1 U14923 ( .ip1(n13672), .ip2(n13671), .op(n13673) );
  inv_1 U14924 ( .ip(n13673), .op(n13674) );
  nor2_1 U14925 ( .ip1(n13675), .ip2(n13674), .op(n13740) );
  inv_1 U14926 ( .ip(n10189), .op(n16838) );
  or2_1 U14927 ( .ip1(n20727), .ip2(n16838), .op(n13677) );
  nor2_1 U14928 ( .ip1(n16423), .ip2(n13676), .op(n13951) );
  inv_1 U14929 ( .ip(n13951), .op(n13847) );
  nand2_1 U14930 ( .ip1(n13677), .ip2(n13847), .op(n13683) );
  or2_1 U14931 ( .ip1(n20220), .ip2(n20221), .op(n13681) );
  inv_1 U14932 ( .ip(n13679), .op(n13680) );
  nand2_1 U14933 ( .ip1(n13681), .ip2(n13680), .op(n13682) );
  nor2_1 U14934 ( .ip1(n13683), .ip2(n13682), .op(n13684) );
  nand2_1 U14935 ( .ip1(n13685), .ip2(n13684), .op(n13687) );
  nor2_1 U14936 ( .ip1(n13687), .ip2(n13686), .op(n13738) );
  inv_1 U14937 ( .ip(n17040), .op(n17043) );
  nand2_1 U14938 ( .ip1(n12932), .ip2(n17043), .op(n13912) );
  inv_1 U14939 ( .ip(n13912), .op(n13689) );
  nor2_1 U14940 ( .ip1(n12932), .ip2(n17043), .op(n13690) );
  nor2_1 U14941 ( .ip1(n13689), .ip2(n13688), .op(n13695) );
  nand2_1 U14942 ( .ip1(n13878), .ip2(n10185), .op(n13693) );
  or2_1 U14943 ( .ip1(n16445), .ip2(n10194), .op(n13692) );
  inv_1 U14944 ( .ip(n13690), .op(n13691) );
  nand2_1 U14945 ( .ip1(n13692), .ip2(n13691), .op(n13718) );
  or2_1 U14946 ( .ip1(n13693), .ip2(n13718), .op(n13694) );
  nand2_1 U14947 ( .ip1(n13695), .ip2(n13694), .op(n13701) );
  inv_1 U14948 ( .ip(n16972), .op(n13708) );
  nor2_1 U14949 ( .ip1(n13708), .ip2(n13707), .op(n13710) );
  inv_1 U14950 ( .ip(n13710), .op(n13697) );
  inv_1 U14951 ( .ip(n17457), .op(n17455) );
  or2_1 U14952 ( .ip1(n17456), .ip2(n17455), .op(n13696) );
  nand2_1 U14953 ( .ip1(n13697), .ip2(n13696), .op(n13706) );
  nand2_1 U14954 ( .ip1(n12596), .ip2(n16811), .op(n13704) );
  or2_1 U14955 ( .ip1(n13022), .ip2(n17006), .op(n13699) );
  nand2_1 U14956 ( .ip1(n13704), .ip2(n13699), .op(n13700) );
  nor2_1 U14957 ( .ip1(n13706), .ip2(n13700), .op(n13720) );
  and2_1 U14958 ( .ip1(n13701), .ip2(n13720), .op(n13716) );
  inv_1 U14959 ( .ip(n12596), .op(n13702) );
  nand2_1 U14960 ( .ip1(n13698), .ip2(n13702), .op(n13918) );
  inv_1 U14961 ( .ip(n13918), .op(n13794) );
  nand2_1 U14962 ( .ip1(n13022), .ip2(n17006), .op(n13917) );
  nor2_1 U14963 ( .ip1(n13794), .ip2(n10229), .op(n13705) );
  or2_1 U14964 ( .ip1(n13706), .ip2(n13705), .op(n13714) );
  inv_1 U14965 ( .ip(n13707), .op(n13877) );
  inv_1 U14966 ( .ip(n13877), .op(n16973) );
  nand2_1 U14967 ( .ip1(n17456), .ip2(n17455), .op(n13711) );
  nor2_1 U14968 ( .ip1(n13711), .ip2(n13710), .op(n13712) );
  nor2_1 U14969 ( .ip1(n13709), .ip2(n13712), .op(n13713) );
  nand2_1 U14970 ( .ip1(n13714), .ip2(n13713), .op(n13715) );
  nor2_1 U14971 ( .ip1(n13716), .ip2(n13715), .op(n13736) );
  nor2_1 U14972 ( .ip1(n13878), .ip2(n13717), .op(n13928) );
  nor2_1 U14973 ( .ip1(n13718), .ip2(n13928), .op(n13719) );
  nand2_1 U14974 ( .ip1(n13720), .ip2(n13719), .op(n13734) );
  inv_1 U14975 ( .ip(n13807), .op(n17480) );
  nand2_1 U14976 ( .ip1(n13808), .ip2(n17479), .op(n13724) );
  nand2_1 U14977 ( .ip1(n13166), .ip2(n17492), .op(n13731) );
  nand2_1 U14978 ( .ip1(n10207), .ip2(n10184), .op(n13810) );
  or2_1 U14979 ( .ip1(n13729), .ip2(n13810), .op(n13730) );
  nand2_1 U14980 ( .ip1(n13731), .ip2(n13730), .op(n13732) );
  nor2_1 U14981 ( .ip1(n13936), .ip2(n13732), .op(n13733) );
  or2_1 U14982 ( .ip1(n13734), .ip2(n13733), .op(n13735) );
  nand2_1 U14983 ( .ip1(n13736), .ip2(n13735), .op(n13737) );
  nand2_1 U14984 ( .ip1(n13738), .ip2(n13737), .op(n13739) );
  nor2_1 U14985 ( .ip1(n13743), .ip2(n13742), .op(n13982) );
  nor2_1 U14986 ( .ip1(n13983), .ip2(n13982), .op(n13744) );
  nand2_1 U14987 ( .ip1(n13744), .ip2(n13977), .op(n13745) );
  nor2_1 U14988 ( .ip1(n13745), .ip2(n13597), .op(n13747) );
  nand3_2 U14989 ( .ip1(n13752), .ip2(n13751), .ip3(n13750), .op(n21531) );
  nor2_1 U14990 ( .ip1(n16479), .ip2(n17819), .op(n17665) );
  nor2_1 U14991 ( .ip1(n13578), .ip2(n13895), .op(n16496) );
  inv_1 U14992 ( .ip(n13755), .op(n13757) );
  inv_1 U14993 ( .ip(n13993), .op(n13759) );
  nand2_1 U14994 ( .ip1(n13854), .ip2(n13855), .op(n13756) );
  nor2_1 U14995 ( .ip1(n13759), .ip2(n13756), .op(n13761) );
  nand2_1 U14996 ( .ip1(n13761), .ip2(n13996), .op(n13790) );
  or2_1 U14997 ( .ip1(n13757), .ip2(n13790), .op(n13764) );
  nand2_1 U14998 ( .ip1(n13906), .ip2(n13758), .op(n13762) );
  inv_1 U14999 ( .ip(n13884), .op(n14007) );
  nor2_1 U15000 ( .ip1(n13759), .ip2(n13615), .op(n13760) );
  not_ab_or_c_or_d U15001 ( .ip1(n13762), .ip2(n13761), .ip3(n14007), .ip4(
        n13760), .op(n13763) );
  nand2_1 U15002 ( .ip1(n13764), .ip2(n13763), .op(n13769) );
  inv_1 U15003 ( .ip(n13981), .op(n13844) );
  nand3_1 U15004 ( .ip1(n13844), .ip2(n13985), .ip3(n13994), .op(n13771) );
  nor2_1 U15005 ( .ip1(n13765), .ip2(n13771), .op(n13767) );
  inv_1 U15006 ( .ip(n13984), .op(n13766) );
  nand3_1 U15007 ( .ip1(n13995), .ip2(n13974), .ip3(n13975), .op(n13777) );
  nand2_1 U15008 ( .ip1(n13767), .ip2(n13775), .op(n13791) );
  inv_1 U15009 ( .ip(n13791), .op(n13768) );
  nand2_1 U15010 ( .ip1(n13769), .ip2(n13768), .op(n13786) );
  inv_1 U15011 ( .ip(n14006), .op(n14014) );
  nand2_1 U15012 ( .ip1(n13902), .ip2(n13985), .op(n13772) );
  inv_1 U15013 ( .ip(n13982), .op(n13861) );
  inv_1 U15014 ( .ip(n13777), .op(n13781) );
  inv_1 U15015 ( .ip(n13904), .op(n13780) );
  nand2_1 U15016 ( .ip1(n13781), .ip2(n13780), .op(n13784) );
  nand2_1 U15017 ( .ip1(n13995), .ip2(n13597), .op(n13782) );
  nand2_1 U15018 ( .ip1(n13786), .ip2(n10203), .op(n13787) );
  inv_1 U15019 ( .ip(n13787), .op(n13842) );
  nand3_1 U15020 ( .ip1(n13997), .ip2(n13885), .ip3(n13956), .op(n13788) );
  or2_1 U15021 ( .ip1(n13788), .ip2(n13961), .op(n13789) );
  or2_1 U15022 ( .ip1(n13790), .ip2(n13789), .op(n13792) );
  nor2_1 U15023 ( .ip1(n13792), .ip2(n13791), .op(n13840) );
  nand3_1 U15024 ( .ip1(n13912), .ip2(n13911), .ip3(n13917), .op(n13819) );
  nor2_1 U15025 ( .ip1(n13913), .ip2(n13819), .op(n13798) );
  inv_1 U15026 ( .ip(n13927), .op(n13793) );
  inv_1 U15027 ( .ip(n13925), .op(n13860) );
  nand3_1 U15028 ( .ip1(n13793), .ip2(n13860), .ip3(n13846), .op(n13828) );
  nor2_1 U15029 ( .ip1(n13794), .ip2(n13828), .op(n13795) );
  nand2_1 U15030 ( .ip1(n13796), .ip2(n13795), .op(n13822) );
  inv_1 U15031 ( .ip(n13822), .op(n13797) );
  nand2_1 U15032 ( .ip1(n13798), .ip2(n13797), .op(n13799) );
  inv_1 U15033 ( .ip(n13799), .op(n13817) );
  nand2_1 U15034 ( .ip1(n19193), .ip2(n13728), .op(n13800) );
  nand2_1 U15035 ( .ip1(n10184), .ip2(n13166), .op(n13802) );
  nand2_1 U15036 ( .ip1(n13881), .ip2(n10207), .op(n18918) );
  inv_1 U15037 ( .ip(n18918), .op(n19427) );
  nand2_1 U15038 ( .ip1(n13802), .ip2(n18918), .op(n13803) );
  or2_1 U15039 ( .ip1(n13801), .ip2(n13803), .op(n13815) );
  inv_1 U15040 ( .ip(n13804), .op(n13805) );
  nand2_1 U15041 ( .ip1(n13805), .ip2(n17480), .op(n13806) );
  nand2_1 U15042 ( .ip1(n13806), .ip2(n17479), .op(n13813) );
  nor2_1 U15043 ( .ip1(n16487), .ip2(n17480), .op(n16507) );
  inv_1 U15044 ( .ip(n17480), .op(n13808) );
  nand2_1 U15045 ( .ip1(n13524), .ip2(n13808), .op(n13809) );
  nand2_1 U15046 ( .ip1(n13810), .ip2(n13809), .op(n13811) );
  not_ab_or_c_or_d U15047 ( .ip1(n13166), .ip2(n17492), .ip3(n16507), .ip4(
        n13811), .op(n13812) );
  nand2_1 U15048 ( .ip1(n13813), .ip2(n13812), .op(n13814) );
  nand2_1 U15049 ( .ip1(n13815), .ip2(n13814), .op(n13816) );
  nand2_1 U15050 ( .ip1(n13817), .ip2(n13816), .op(n13838) );
  inv_1 U15051 ( .ip(n13933), .op(n13818) );
  nor2_1 U15052 ( .ip1(n13818), .ip2(n13928), .op(n13820) );
  nor2_1 U15053 ( .ip1(n13820), .ip2(n13819), .op(n13821) );
  not_ab_or_c_or_d U15054 ( .ip1(n13914), .ip2(n13917), .ip3(n13915), .ip4(
        n13821), .op(n13823) );
  nor2_1 U15055 ( .ip1(n13823), .ip2(n13822), .op(n13836) );
  inv_1 U15056 ( .ip(n13924), .op(n13824) );
  nand2_1 U15057 ( .ip1(n13846), .ip2(n13824), .op(n13825) );
  nand2_1 U15058 ( .ip1(n13825), .ip2(n13847), .op(n13830) );
  inv_1 U15059 ( .ip(n13921), .op(n13826) );
  nor2_1 U15060 ( .ip1(n13557), .ip2(n13826), .op(n13827) );
  nor2_1 U15061 ( .ip1(n13828), .ip2(n13827), .op(n13829) );
  nor2_1 U15062 ( .ip1(n13830), .ip2(n13829), .op(n13831) );
  or2_1 U15063 ( .ip1(n13832), .ip2(n13831), .op(n13834) );
  nand2_1 U15064 ( .ip1(n13834), .ip2(n13833), .op(n13835) );
  nor2_1 U15065 ( .ip1(n13836), .ip2(n13835), .op(n13837) );
  nand2_1 U15066 ( .ip1(n13838), .ip2(n13837), .op(n13839) );
  nand2_1 U15067 ( .ip1(n13840), .ip2(n13839), .op(n13841) );
  nand2_1 U15068 ( .ip1(n13842), .ip2(n13841), .op(n13843) );
  nand2_1 U15069 ( .ip1(n13845), .ip2(n13844), .op(n16932) );
  nand2_1 U15070 ( .ip1(n13954), .ip2(n13956), .op(n16858) );
  nand2_1 U15071 ( .ip1(n13899), .ip2(n13974), .op(n17099) );
  nand2_1 U15072 ( .ip1(n13960), .ip2(n13963), .op(n19438) );
  nand2_1 U15073 ( .ip1(n13847), .ip2(n13846), .op(n16688) );
  nand2_1 U15074 ( .ip1(n13930), .ip2(n13912), .op(n17046) );
  nand2_1 U15075 ( .ip1(n13933), .ip2(n13911), .op(n17588) );
  nand2_1 U15076 ( .ip1(n13995), .ip2(n13900), .op(n20910) );
  nand2_1 U15077 ( .ip1(n13615), .ip2(n13854), .op(n17177) );
  nand2_1 U15078 ( .ip1(n13758), .ip2(n13855), .op(n17534) );
  nand2_1 U15079 ( .ip1(n13921), .ip2(n13860), .op(n17461) );
  nand2_1 U15080 ( .ip1(n13861), .ip2(n13985), .op(n19203) );
  nand2_1 U15081 ( .ip1(n13863), .ip2(n13862), .op(n20226) );
  nor2_2 U15082 ( .ip1(n13867), .ip2(n13866), .op(n13893) );
  xor2_1 U15083 ( .ip1(n20727), .ip2(n13627), .op(n20729) );
  xnor2_1 U15084 ( .ip1(n16418), .ip2(n13868), .op(n16494) );
  xnor2_1 U15085 ( .ip1(n13698), .ip2(n12596), .op(n16809) );
  xor2_1 U15086 ( .ip1(n10198), .ip2(n10184), .op(n16717) );
  inv_1 U15087 ( .ip(n16717), .op(n13872) );
  xnor2_1 U15088 ( .ip1(n16487), .ip2(n13524), .op(n13871) );
  nand2_1 U15089 ( .ip1(n16809), .ip2(n13873), .op(n13874) );
  inv_1 U15090 ( .ip(n13874), .op(n13875) );
  xor2_1 U15091 ( .ip1(n10186), .ip2(n18731), .op(n18735) );
  xnor2_1 U15092 ( .ip1(n16972), .ip2(n13877), .op(n16970) );
  xor2_1 U15093 ( .ip1(n17480), .ip2(n17479), .op(n17483) );
  nor2_1 U15094 ( .ip1(n16970), .ip2(n17483), .op(n13879) );
  nand2_1 U15095 ( .ip1(n13879), .ip2(n10177), .op(n13880) );
  nor2_1 U15096 ( .ip1(n18735), .ip2(n13880), .op(n13883) );
  inv_1 U15097 ( .ip(n11180), .op(n17270) );
  xor2_1 U15098 ( .ip1(n17277), .ip2(n17270), .op(n17280) );
  xor2_1 U15099 ( .ip1(n13881), .ip2(n17492), .op(n16754) );
  nand2_1 U15100 ( .ip1(n13993), .ip2(n13884), .op(n16598) );
  nand2_1 U15101 ( .ip1(n13886), .ip2(n13885), .op(n16637) );
  inv_1 U15102 ( .ip(n13887), .op(n13888) );
  nand2_1 U15103 ( .ip1(n13889), .ip2(n13888), .op(n17141) );
  nand2_1 U15104 ( .ip1(n13932), .ip2(n13917), .op(n17010) );
  nand2_2 U15105 ( .ip1(n13893), .ip2(n13892), .op(n13897) );
  nand2_1 U15106 ( .ip1(n13897), .ip2(n13894), .op(n14023) );
  inv_1 U15107 ( .ip(n13895), .op(n13896) );
  or2_1 U15108 ( .ip1(n13578), .ip2(n13896), .op(n16485) );
  nor2_2 U15109 ( .ip1(n16485), .ip2(n13897), .op(n13898) );
  nor2_2 U15110 ( .ip1(n16913), .ip2(n13898), .op(n14022) );
  nand2_1 U15111 ( .ip1(n13905), .ip2(n13995), .op(n13991) );
  inv_1 U15112 ( .ip(n13906), .op(n14000) );
  or2_1 U15113 ( .ip1(n14000), .ip2(n14001), .op(n13907) );
  nor4_1 U15114 ( .ip1(n14007), .ip2(n13908), .ip3(n14006), .ip4(n13907), .op(
        n13909) );
  nand2_1 U15115 ( .ip1(n13933), .ip2(n13913), .op(n13916) );
  inv_1 U15116 ( .ip(n13930), .op(n13914) );
  ab_or_c_or_d U15117 ( .ip1(n10228), .ip2(n13916), .ip3(n13915), .ip4(n13914), 
        .op(n13920) );
  nand2_1 U15118 ( .ip1(n13920), .ip2(n13919), .op(n13923) );
  nand2_1 U15119 ( .ip1(n13923), .ip2(n13935), .op(n13946) );
  nor2_1 U15120 ( .ip1(n13927), .ip2(n13926), .op(n13945) );
  inv_1 U15121 ( .ip(n13928), .op(n13929) );
  inv_1 U15122 ( .ip(n18918), .op(n16670) );
  nand2_1 U15123 ( .ip1(n16670), .ip2(n10184), .op(n13938) );
  nand2_1 U15124 ( .ip1(n13938), .ip2(n10195), .op(n13939) );
  nand2_1 U15125 ( .ip1(n10226), .ip2(n13943), .op(n13944) );
  nand3_1 U15126 ( .ip1(n13946), .ip2(n13945), .ip3(n13944), .op(n13953) );
  nor2_1 U15127 ( .ip1(n13948), .ip2(n13947), .op(n13949) );
  nand2_1 U15128 ( .ip1(n13949), .ip2(n13954), .op(n13958) );
  nor4_1 U15129 ( .ip1(n12139), .ip2(n13951), .ip3(n13950), .ip4(n13958), .op(
        n13952) );
  nand2_1 U15130 ( .ip1(n13953), .ip2(n13952), .op(n13972) );
  nand2_1 U15131 ( .ip1(n13955), .ip2(n13954), .op(n13957) );
  nand2_1 U15132 ( .ip1(n13957), .ip2(n13956), .op(n13970) );
  nor2_1 U15133 ( .ip1(n13970), .ip2(n13969), .op(n13971) );
  nand2_1 U15134 ( .ip1(n13972), .ip2(n13971), .op(n13973) );
  nand2_1 U15135 ( .ip1(n13910), .ip2(n13973), .op(n14019) );
  nor2_1 U15136 ( .ip1(n13597), .ip2(n13978), .op(n13979) );
  or3_1 U15137 ( .ip1(n13983), .ip2(n13982), .ip3(n13844), .op(n13988) );
  nand2_1 U15138 ( .ip1(n13985), .ip2(n13984), .op(n13986) );
  nand2_1 U15139 ( .ip1(n13986), .ip2(n13779), .op(n13987) );
  inv_1 U15140 ( .ip(n13991), .op(n14016) );
  nand2_1 U15141 ( .ip1(n13993), .ip2(n13992), .op(n14013) );
  nand2_1 U15142 ( .ip1(n13995), .ip2(n13994), .op(n14012) );
  nand2_1 U15143 ( .ip1(n13997), .ip2(n13996), .op(n13998) );
  inv_1 U15144 ( .ip(n13998), .op(n13999) );
  nor2_1 U15145 ( .ip1(n14000), .ip2(n13999), .op(n14003) );
  inv_1 U15146 ( .ip(n14001), .op(n14002) );
  nand2_1 U15147 ( .ip1(n14003), .ip2(n14002), .op(n14004) );
  nand2_1 U15148 ( .ip1(n14005), .ip2(n14004), .op(n14009) );
  nor2_1 U15149 ( .ip1(n14007), .ip2(n14006), .op(n14008) );
  nand2_1 U15150 ( .ip1(n14009), .ip2(n14008), .op(n14010) );
  inv_1 U15151 ( .ip(n14010), .op(n14011) );
  not_ab_or_c_or_d U15152 ( .ip1(n14014), .ip2(n14013), .ip3(n14012), .ip4(
        n14011), .op(n14015) );
  nor2_1 U15153 ( .ip1(n14016), .ip2(n14015), .op(n14017) );
  nor2_1 U15154 ( .ip1(n13990), .ip2(n14017), .op(n14018) );
  nand4_2 U15155 ( .ip1(n14024), .ip2(n14023), .ip3(n14022), .ip4(n14021), 
        .op(n17666) );
  nand2_4 U15156 ( .ip1(n10211), .ip2(n17666), .op(n14129) );
  nand2_4 U15157 ( .ip1(n14392), .ip2(n14129), .op(n14074) );
  inv_1 U15158 ( .ip(n17779), .op(n14027) );
  inv_1 U15159 ( .ip(n14025), .op(n14026) );
  nor2_1 U15160 ( .ip1(n14027), .ip2(n14026), .op(n14028) );
  nand2_1 U15161 ( .ip1(n17891), .ip2(n14028), .op(n21088) );
  inv_1 U15162 ( .ip(n17888), .op(n14167) );
  and2_1 U15163 ( .ip1(n21088), .ip2(n14167), .op(n17669) );
  inv_1 U15164 ( .ip(n14090), .op(n14310) );
  nand2_1 U15165 ( .ip1(n14340), .ip2(\pipeline/PC_DX [24]), .op(n14041) );
  inv_1 U15166 ( .ip(n17669), .op(n14033) );
  nand2_1 U15167 ( .ip1(n14033), .ip2(n14032), .op(n14035) );
  nand2_2 U15168 ( .ip1(n10238), .ip2(n14129), .op(n14157) );
  inv_2 U15169 ( .ip(n14157), .op(n14080) );
  inv_1 U15170 ( .ip(n20611), .op(n16112) );
  nor2_1 U15171 ( .ip1(n16112), .ip2(n14392), .op(n14039) );
  inv_1 U15172 ( .ip(n21088), .op(n20975) );
  and2_1 U15173 ( .ip1(n14169), .ip2(n20975), .op(n14466) );
  nand2_1 U15174 ( .ip1(n14466), .ip2(\pipeline/epc [24]), .op(n14037) );
  nand2_1 U15175 ( .ip1(n10364), .ip2(\pipeline/csr/mtvec [24]), .op(n14036)
         );
  nand2_1 U15176 ( .ip1(n14037), .ip2(n14036), .op(n14038) );
  not_ab_or_c_or_d U15177 ( .ip1(\pipeline/PC_IF [24]), .ip2(n14404), .ip3(
        n14039), .ip4(n14038), .op(n14040) );
  inv_1 U15178 ( .ip(n15401), .op(n20278) );
  nor2_1 U15179 ( .ip1(n20278), .ip2(n14392), .op(n14045) );
  nand2_1 U15180 ( .ip1(n14466), .ip2(\pipeline/epc [23]), .op(n14043) );
  nand2_1 U15181 ( .ip1(n10364), .ip2(\pipeline/csr/mtvec [23]), .op(n14042)
         );
  nand2_1 U15182 ( .ip1(n14043), .ip2(n14042), .op(n14044) );
  not_ab_or_c_or_d U15183 ( .ip1(\pipeline/PC_IF [23]), .ip2(n14404), .ip3(
        n14045), .ip4(n14044), .op(n14047) );
  nand2_1 U15184 ( .ip1(n18021), .ip2(\pipeline/PC_DX [23]), .op(n14046) );
  nor2_1 U15185 ( .ip1(n14497), .ip2(n14503), .op(n14049) );
  inv_1 U15186 ( .ip(n14435), .op(n14048) );
  nor2_1 U15187 ( .ip1(n14049), .ip2(n14048), .op(n14390) );
  nand2_1 U15188 ( .ip1(\pipeline/PC_DX [21]), .ip2(n14413), .op(n14055) );
  inv_1 U15189 ( .ip(n20586), .op(n15531) );
  nor2_1 U15190 ( .ip1(n15531), .ip2(n14392), .op(n14053) );
  nand2_1 U15191 ( .ip1(n14466), .ip2(\pipeline/epc [21]), .op(n14051) );
  nand2_1 U15192 ( .ip1(n10364), .ip2(\pipeline/csr/mtvec [21]), .op(n14050)
         );
  nand2_1 U15193 ( .ip1(n14051), .ip2(n14050), .op(n14052) );
  not_ab_or_c_or_d U15194 ( .ip1(\pipeline/PC_IF [21]), .ip2(n14404), .ip3(
        n14053), .ip4(n14052), .op(n14054) );
  inv_2 U15195 ( .ip(n14235), .op(n14399) );
  nand2_1 U15196 ( .ip1(n14399), .ip2(\pipeline/PC_DX [22]), .op(n14065) );
  nand2_1 U15197 ( .ip1(n14057), .ip2(n14056), .op(n14058) );
  nand2_1 U15198 ( .ip1(n14059), .ip2(n14058), .op(n15369) );
  inv_1 U15199 ( .ip(n15369), .op(n20599) );
  nor2_1 U15200 ( .ip1(n20599), .ip2(n14392), .op(n14063) );
  nand2_1 U15201 ( .ip1(n14466), .ip2(\pipeline/epc [22]), .op(n14061) );
  nand2_1 U15202 ( .ip1(n10364), .ip2(\pipeline/csr/mtvec [22]), .op(n14060)
         );
  nand2_1 U15203 ( .ip1(n14061), .ip2(n14060), .op(n14062) );
  not_ab_or_c_or_d U15204 ( .ip1(\pipeline/PC_IF [22]), .ip2(n14404), .ip3(
        n14063), .ip4(n14062), .op(n14064) );
  mux2_1 U15205 ( .ip1(n14503), .ip2(n14511), .s(n14504), .op(n14436) );
  inv_1 U15206 ( .ip(n15693), .op(n20424) );
  nor2_1 U15207 ( .ip1(n20424), .ip2(n14392), .op(n14069) );
  nand2_1 U15208 ( .ip1(n14466), .ip2(\pipeline/epc [14]), .op(n14067) );
  nand2_1 U15209 ( .ip1(n10364), .ip2(\pipeline/csr/mtvec [14]), .op(n14066)
         );
  nand2_1 U15210 ( .ip1(n14067), .ip2(n14066), .op(n14068) );
  nand2_1 U15211 ( .ip1(n14073), .ip2(n14072), .op(n14120) );
  inv_1 U15212 ( .ip(n14120), .op(n14077) );
  nand2_1 U15213 ( .ip1(n14031), .ip2(\pipeline/dmem_type[2] ), .op(n14075) );
  inv_1 U15214 ( .ip(n14074), .op(n14243) );
  nand2_1 U15215 ( .ip1(n14075), .ip2(n14337), .op(n14119) );
  nand2_1 U15216 ( .ip1(\pipeline/PC_DX [13]), .ip2(n14399), .op(n14086) );
  inv_1 U15217 ( .ip(n20400), .op(n15467) );
  nor2_1 U15218 ( .ip1(n15467), .ip2(n14392), .op(n14084) );
  nand2_1 U15219 ( .ip1(n14466), .ip2(\pipeline/epc [13]), .op(n14082) );
  nand2_1 U15220 ( .ip1(n10364), .ip2(\pipeline/csr/mtvec [13]), .op(n14081)
         );
  nand2_1 U15221 ( .ip1(n14082), .ip2(n14081), .op(n14083) );
  not_ab_or_c_or_d U15222 ( .ip1(\pipeline/PC_IF [13]), .ip2(n18024), .ip3(
        n14084), .ip4(n14083), .op(n14085) );
  nand2_1 U15223 ( .ip1(n14086), .ip2(n14085), .op(n14223) );
  nand2_1 U15224 ( .ip1(n14031), .ip2(dmem_hsize[1]), .op(n14087) );
  and2_1 U15225 ( .ip1(n14087), .ip2(n14337), .op(n14224) );
  inv_1 U15226 ( .ip(n14224), .op(n14088) );
  nand2_1 U15227 ( .ip1(n14223), .ip2(n14088), .op(n14364) );
  nand2_1 U15228 ( .ip1(n14031), .ip2(\pipeline/inst_DX [17]), .op(n14089) );
  inv_1 U15229 ( .ip(\pipeline/PC_DX [17]), .op(n14091) );
  or2_1 U15230 ( .ip1(n14339), .ip2(n14091), .op(n14097) );
  inv_1 U15231 ( .ip(n20007), .op(n15499) );
  nor2_1 U15232 ( .ip1(n15499), .ip2(n14392), .op(n14095) );
  nand2_1 U15233 ( .ip1(n14466), .ip2(\pipeline/epc [17]), .op(n14093) );
  nand2_1 U15234 ( .ip1(n10364), .ip2(\pipeline/csr/mtvec [17]), .op(n14092)
         );
  nand2_1 U15235 ( .ip1(n14093), .ip2(n14092), .op(n14094) );
  not_ab_or_c_or_d U15236 ( .ip1(\pipeline/PC_IF [17]), .ip2(n14404), .ip3(
        n14095), .ip4(n14094), .op(n14096) );
  nand2_1 U15237 ( .ip1(n14097), .ip2(n14096), .op(n14348) );
  xnor2_1 U15238 ( .ip1(n14349), .ip2(n14348), .op(n14361) );
  inv_1 U15239 ( .ip(\pipeline/PC_DX [16]), .op(n14098) );
  or2_1 U15240 ( .ip1(n14098), .ip2(n14310), .op(n14104) );
  inv_1 U15241 ( .ip(n14593), .op(n18148) );
  nor2_1 U15242 ( .ip1(n18148), .ip2(n14392), .op(n14102) );
  nand2_1 U15243 ( .ip1(n14466), .ip2(\pipeline/epc [16]), .op(n14100) );
  nand2_1 U15244 ( .ip1(n10364), .ip2(\pipeline/csr/mtvec [16]), .op(n14099)
         );
  nand2_1 U15245 ( .ip1(n14100), .ip2(n14099), .op(n14101) );
  not_ab_or_c_or_d U15246 ( .ip1(\pipeline/PC_IF [16]), .ip2(n14404), .ip3(
        n14102), .ip4(n14101), .op(n14103) );
  nand2_1 U15247 ( .ip1(n14104), .ip2(n14103), .op(n14107) );
  nand2_1 U15248 ( .ip1(n14031), .ip2(\pipeline/inst_DX [16]), .op(n14105) );
  and2_1 U15249 ( .ip1(n14105), .ip2(n14337), .op(n14108) );
  inv_1 U15250 ( .ip(n14108), .op(n14106) );
  nand2_1 U15251 ( .ip1(n14107), .ip2(n14106), .op(n14362) );
  nand2_1 U15252 ( .ip1(n14361), .ip2(n14362), .op(n14440) );
  xnor2_1 U15253 ( .ip1(n14108), .ip2(n14107), .op(n14371) );
  inv_1 U15254 ( .ip(n20426), .op(n15726) );
  nor2_1 U15255 ( .ip1(n15726), .ip2(n14392), .op(n14112) );
  nand2_1 U15256 ( .ip1(n14466), .ip2(\pipeline/epc [15]), .op(n14110) );
  nand2_1 U15257 ( .ip1(n10364), .ip2(\pipeline/csr/mtvec [15]), .op(n14109)
         );
  nand2_1 U15258 ( .ip1(n14110), .ip2(n14109), .op(n14111) );
  not_ab_or_c_or_d U15259 ( .ip1(\pipeline/PC_IF [15]), .ip2(n18024), .ip3(
        n14112), .ip4(n14111), .op(n14113) );
  nand2_1 U15260 ( .ip1(n14031), .ip2(\pipeline/inst_DX [15]), .op(n14115) );
  nand2_1 U15261 ( .ip1(n14115), .ip2(n14337), .op(n14117) );
  nand2_1 U15262 ( .ip1(n14118), .ip2(n14117), .op(n14373) );
  inv_1 U15263 ( .ip(n14373), .op(n14116) );
  or2_1 U15264 ( .ip1(n14371), .ip2(n14116), .op(n18285) );
  xnor2_1 U15265 ( .ip1(n14117), .ip2(n14118), .op(n14366) );
  nand2_1 U15266 ( .ip1(n14120), .ip2(n14119), .op(n14367) );
  inv_1 U15267 ( .ip(n14438), .op(n14309) );
  nand2_1 U15268 ( .ip1(\pipeline/PC_DX [8]), .ip2(n14413), .op(n14128) );
  nand2_1 U15269 ( .ip1(n14122), .ip2(n14121), .op(n15433) );
  nor2_1 U15270 ( .ip1(n15433), .ip2(n14392), .op(n14126) );
  nand2_1 U15271 ( .ip1(n14466), .ip2(\pipeline/epc [8]), .op(n14124) );
  nand2_1 U15272 ( .ip1(n10364), .ip2(\pipeline/csr/mtvec [8]), .op(n14123) );
  nand2_1 U15273 ( .ip1(n14124), .ip2(n14123), .op(n14125) );
  not_ab_or_c_or_d U15274 ( .ip1(\pipeline/PC_IF [8]), .ip2(n18024), .ip3(
        n14126), .ip4(n14125), .op(n14127) );
  nand2_1 U15275 ( .ip1(n14128), .ip2(n14127), .op(n14265) );
  nand2_1 U15276 ( .ip1(n14129), .ip2(n14029), .op(n14318) );
  and2_1 U15277 ( .ip1(n14318), .ip2(\pipeline/inst_DX [28]), .op(n14266) );
  and2_1 U15278 ( .ip1(n14265), .ip2(n14266), .op(n19688) );
  inv_1 U15279 ( .ip(n20485), .op(n15962) );
  nor2_1 U15280 ( .ip1(n15962), .ip2(n14392), .op(n14133) );
  nand2_1 U15281 ( .ip1(n14466), .ip2(\pipeline/epc [6]), .op(n14131) );
  nand2_1 U15282 ( .ip1(n10364), .ip2(\pipeline/prv [1]), .op(n14130) );
  nand2_1 U15283 ( .ip1(n14131), .ip2(n14130), .op(n14132) );
  not_ab_or_c_or_d U15284 ( .ip1(\pipeline/PC_IF [6]), .ip2(n18024), .ip3(
        n14133), .ip4(n14132), .op(n14135) );
  nand2_1 U15285 ( .ip1(\pipeline/PC_DX [6]), .ip2(n14399), .op(n14134) );
  nand2_1 U15286 ( .ip1(n14135), .ip2(n14134), .op(n14217) );
  nand2_1 U15287 ( .ip1(n14318), .ip2(\pipeline/inst_DX [26]), .op(n14137) );
  nand2_1 U15288 ( .ip1(n10364), .ip2(\pipeline/csr/mtvec [6]), .op(n14136) );
  nand2_1 U15289 ( .ip1(n14137), .ip2(n14136), .op(n14218) );
  and2_1 U15290 ( .ip1(n14217), .ip2(n14218), .op(n18232) );
  nand2_1 U15291 ( .ip1(n14413), .ip2(\pipeline/PC_DX [7]), .op(n14143) );
  inv_1 U15292 ( .ip(n15928), .op(n20381) );
  nor2_1 U15293 ( .ip1(n20381), .ip2(n14392), .op(n14141) );
  nand2_1 U15294 ( .ip1(n14466), .ip2(\pipeline/epc [7]), .op(n14139) );
  nand2_1 U15295 ( .ip1(n10364), .ip2(\pipeline/csr/mtvec [7]), .op(n14138) );
  nand2_1 U15296 ( .ip1(n14139), .ip2(n14138), .op(n14140) );
  not_ab_or_c_or_d U15297 ( .ip1(\pipeline/PC_IF [7]), .ip2(n18024), .ip3(
        n14141), .ip4(n14140), .op(n14142) );
  nand2_1 U15298 ( .ip1(n14143), .ip2(n14142), .op(n14146) );
  inv_1 U15299 ( .ip(n14146), .op(n14145) );
  and2_1 U15300 ( .ip1(n14318), .ip2(\pipeline/inst_DX [27]), .op(n14147) );
  inv_1 U15301 ( .ip(n14147), .op(n14144) );
  nand2_1 U15302 ( .ip1(n14145), .ip2(n14144), .op(n18228) );
  nand2_1 U15303 ( .ip1(n18232), .ip2(n18228), .op(n14148) );
  nand2_1 U15304 ( .ip1(n14147), .ip2(n14146), .op(n18227) );
  nand2_1 U15305 ( .ip1(n14148), .ip2(n18227), .op(n14580) );
  nor2_1 U15306 ( .ip1(n19688), .ip2(n14580), .op(n14222) );
  nand2_1 U15307 ( .ip1(n14090), .ip2(\pipeline/PC_DX [2]), .op(n14156) );
  nand2_1 U15308 ( .ip1(n14466), .ip2(\pipeline/epc [2]), .op(n14150) );
  nand2_1 U15309 ( .ip1(n10364), .ip2(\pipeline/csr/mtvec [2]), .op(n14149) );
  nand2_1 U15310 ( .ip1(n14150), .ip2(n14149), .op(n14152) );
  inv_1 U15311 ( .ip(n15789), .op(n17345) );
  nor2_1 U15312 ( .ip1(n17345), .ip2(n14392), .op(n14151) );
  nor2_1 U15313 ( .ip1(n14152), .ip2(n14151), .op(n14154) );
  nand2_1 U15314 ( .ip1(\pipeline/PC_IF [2]), .ip2(n14404), .op(n14153) );
  nand2_1 U15315 ( .ip1(n14156), .ip2(n14155), .op(n17435) );
  nand2_1 U15316 ( .ip1(n14340), .ip2(\pipeline/PC_DX [1]), .op(n14162) );
  inv_1 U15317 ( .ip(n14597), .op(n17334) );
  nor2_1 U15318 ( .ip1(n17334), .ip2(n14392), .op(n14160) );
  inv_1 U15319 ( .ip(\pipeline/PC_IF [1]), .op(n14158) );
  nor2_1 U15320 ( .ip1(n14158), .ip2(n14157), .op(n14159) );
  nor2_1 U15321 ( .ip1(n14160), .ip2(n14159), .op(n14161) );
  inv_1 U15322 ( .ip(n14240), .op(n14186) );
  nand2_1 U15323 ( .ip1(n14186), .ip2(\pipeline/inst_DX [8]), .op(n14164) );
  nand2_1 U15324 ( .ip1(n14241), .ip2(\pipeline/inst_DX [21]), .op(n14163) );
  nand2_1 U15325 ( .ip1(n14164), .ip2(n14163), .op(n21992) );
  inv_1 U15326 ( .ip(\pipeline/inst_DX [9]), .op(n14166) );
  mux2_1 U15327 ( .ip1(\pipeline/inst_DX [22]), .ip2(n14168), .s(n14167), .op(
        n14172) );
  inv_1 U15328 ( .ip(n14169), .op(n14170) );
  nor2_1 U15329 ( .ip1(n20975), .ip2(n14170), .op(n14171) );
  and2_1 U15330 ( .ip1(n14172), .ip2(n14171), .op(n17436) );
  inv_1 U15331 ( .ip(n17436), .op(n14173) );
  nand2_1 U15332 ( .ip1(n17437), .ip2(n14173), .op(n14174) );
  nand2_1 U15333 ( .ip1(n17435), .ip2(n14174), .op(n14176) );
  or2_1 U15334 ( .ip1(n17437), .ip2(n14173), .op(n14175) );
  nand2_2 U15335 ( .ip1(n14176), .ip2(n14175), .op(n21162) );
  nand2_1 U15336 ( .ip1(n14186), .ip2(\pipeline/inst_DX [10]), .op(n14178) );
  nand2_1 U15337 ( .ip1(n14241), .ip2(\pipeline/inst_DX [23]), .op(n14177) );
  nand2_1 U15338 ( .ip1(n14178), .ip2(n14177), .op(n14206) );
  inv_1 U15339 ( .ip(\pipeline/PC_DX [3]), .op(n14179) );
  or2_1 U15340 ( .ip1(n14235), .ip2(n14179), .op(n14185) );
  inv_1 U15341 ( .ip(n15796), .op(n17855) );
  nor2_1 U15342 ( .ip1(n17855), .ip2(n14392), .op(n14183) );
  nand2_1 U15343 ( .ip1(n14466), .ip2(\pipeline/epc [3]), .op(n14181) );
  nand2_1 U15344 ( .ip1(n10364), .ip2(\pipeline/csr/mtvec [3]), .op(n14180) );
  nand2_1 U15345 ( .ip1(n14181), .ip2(n14180), .op(n14182) );
  not_ab_or_c_or_d U15346 ( .ip1(\pipeline/PC_IF [3]), .ip2(n18024), .ip3(
        n14183), .ip4(n14182), .op(n14184) );
  nand2_1 U15347 ( .ip1(n14185), .ip2(n14184), .op(n14207) );
  nor2_1 U15348 ( .ip1(n14206), .ip2(n14207), .op(n21161) );
  nand2_1 U15349 ( .ip1(n14340), .ip2(\pipeline/PC_DX [4]), .op(n14211) );
  nand2_1 U15350 ( .ip1(n14186), .ip2(\pipeline/inst_DX [11]), .op(n14188) );
  nand2_1 U15351 ( .ip1(n14241), .ip2(\pipeline/inst_DX [24]), .op(n14187) );
  nand2_1 U15352 ( .ip1(n14188), .ip2(n14187), .op(n17957) );
  inv_1 U15353 ( .ip(n17957), .op(n14195) );
  inv_1 U15354 ( .ip(n17939), .op(n15661) );
  nor2_1 U15355 ( .ip1(n15661), .ip2(n14392), .op(n14192) );
  nand2_1 U15356 ( .ip1(n14466), .ip2(\pipeline/epc [4]), .op(n14190) );
  nand2_1 U15357 ( .ip1(n10364), .ip2(\pipeline/csr/mtvec [4]), .op(n14189) );
  nand2_1 U15358 ( .ip1(n14190), .ip2(n14189), .op(n14191) );
  inv_1 U15359 ( .ip(n14209), .op(n14196) );
  nand2_2 U15360 ( .ip1(n21162), .ip2(n14197), .op(n17989) );
  inv_1 U15361 ( .ip(n14235), .op(n18021) );
  nand2_1 U15362 ( .ip1(n18021), .ip2(\pipeline/PC_DX [5]), .op(n14203) );
  inv_1 U15363 ( .ip(n20476), .op(n15862) );
  nor2_1 U15364 ( .ip1(n15862), .ip2(n14392), .op(n14201) );
  nand2_1 U15365 ( .ip1(n14466), .ip2(\pipeline/epc [5]), .op(n14199) );
  nand2_1 U15366 ( .ip1(n10364), .ip2(\pipeline/prv [0]), .op(n14198) );
  nand2_1 U15367 ( .ip1(n14199), .ip2(n14198), .op(n14200) );
  not_ab_or_c_or_d U15368 ( .ip1(\pipeline/PC_IF [5]), .ip2(n18024), .ip3(
        n14201), .ip4(n14200), .op(n14202) );
  nand2_1 U15369 ( .ip1(n14203), .ip2(n14202), .op(n14215) );
  nand2_1 U15370 ( .ip1(n14318), .ip2(\pipeline/inst_DX [25]), .op(n14205) );
  nand2_1 U15371 ( .ip1(n10364), .ip2(\pipeline/csr/mtvec [5]), .op(n14204) );
  nand2_1 U15372 ( .ip1(n14205), .ip2(n14204), .op(n14216) );
  and2_1 U15373 ( .ip1(n14215), .ip2(n14216), .op(n21035) );
  nand2_1 U15374 ( .ip1(n14207), .ip2(n14206), .op(n14208) );
  inv_1 U15375 ( .ip(n14208), .op(n21160) );
  nand2_1 U15376 ( .ip1(n21160), .ip2(n14209), .op(n14213) );
  nand2_1 U15377 ( .ip1(n14211), .ip2(n14210), .op(n17956) );
  nand2_1 U15378 ( .ip1(n17956), .ip2(n17957), .op(n14212) );
  nor2_1 U15379 ( .ip1(n14216), .ip2(n14215), .op(n21036) );
  inv_1 U15380 ( .ip(n18228), .op(n14219) );
  nor2_1 U15381 ( .ip1(n14218), .ip2(n14217), .op(n18229) );
  nor3_1 U15382 ( .ip1(n21036), .ip2(n14219), .ip3(n18229), .op(n14220) );
  nand2_1 U15383 ( .ip1(\pipeline/PC_DX [12]), .ip2(n14340), .op(n14231) );
  inv_1 U15384 ( .ip(n16402), .op(n20392) );
  nor2_1 U15385 ( .ip1(n20392), .ip2(n14392), .op(n14229) );
  nand2_1 U15386 ( .ip1(n14466), .ip2(\pipeline/epc [12]), .op(n14227) );
  nand2_1 U15387 ( .ip1(n10364), .ip2(\pipeline/csr/mtvec [12]), .op(n14226)
         );
  nand2_1 U15388 ( .ip1(n14227), .ip2(n14226), .op(n14228) );
  not_ab_or_c_or_d U15389 ( .ip1(\pipeline/PC_IF [12]), .ip2(n18024), .ip3(
        n14229), .ip4(n14228), .op(n14230) );
  nand2_1 U15390 ( .ip1(n14231), .ip2(n14230), .op(n14234) );
  nand2_1 U15391 ( .ip1(n14031), .ip2(dmem_hsize[0]), .op(n14232) );
  nand2_1 U15392 ( .ip1(n14232), .ip2(n14337), .op(n14233) );
  nand2_1 U15393 ( .ip1(n14234), .ip2(n14233), .op(n14303) );
  inv_1 U15394 ( .ip(\pipeline/PC_DX [11]), .op(n14236) );
  or2_1 U15395 ( .ip1(n14236), .ip2(n14235), .op(n14272) );
  inv_1 U15396 ( .ip(n14392), .op(n18023) );
  nand2_1 U15397 ( .ip1(n18023), .ip2(n16226), .op(n14238) );
  nand2_1 U15398 ( .ip1(n14466), .ip2(\pipeline/epc [11]), .op(n14237) );
  and2_1 U15399 ( .ip1(n14238), .ip2(n14237), .op(n14275) );
  nand2_1 U15400 ( .ip1(n14272), .ip2(n14275), .op(n14271) );
  inv_1 U15401 ( .ip(\pipeline/inst_DX [7]), .op(n14239) );
  nor2_1 U15402 ( .ip1(n14240), .ip2(n14239), .op(n14247) );
  nand2_1 U15403 ( .ip1(n14243), .ip2(n14242), .op(n14245) );
  or2_1 U15404 ( .ip1(n15324), .ip2(n14392), .op(n14244) );
  nand2_1 U15405 ( .ip1(n14245), .ip2(n14244), .op(n14246) );
  or2_1 U15406 ( .ip1(n14247), .ip2(n14246), .op(n14276) );
  nand2_1 U15407 ( .ip1(n14271), .ip2(n14276), .op(n14300) );
  and2_1 U15408 ( .ip1(n14318), .ip2(\pipeline/inst_DX [30]), .op(n14285) );
  nand2_1 U15409 ( .ip1(n14413), .ip2(\pipeline/PC_DX [10]), .op(n14255) );
  inv_1 U15410 ( .ip(n14601), .op(n14249) );
  nor2_1 U15411 ( .ip1(n14249), .ip2(n14392), .op(n14253) );
  nand2_1 U15412 ( .ip1(n14466), .ip2(\pipeline/epc [10]), .op(n14251) );
  nand2_1 U15413 ( .ip1(n10364), .ip2(\pipeline/csr/mtvec [10]), .op(n14250)
         );
  nand2_1 U15414 ( .ip1(n14251), .ip2(n14250), .op(n14252) );
  not_ab_or_c_or_d U15415 ( .ip1(\pipeline/PC_IF [10]), .ip2(n18024), .ip3(
        n14253), .ip4(n14252), .op(n14254) );
  nand2_1 U15416 ( .ip1(n14255), .ip2(n14254), .op(n14290) );
  xnor2_1 U15417 ( .ip1(n14285), .ip2(n14290), .op(n14262) );
  and2_1 U15418 ( .ip1(n14318), .ip2(\pipeline/inst_DX [29]), .op(n14264) );
  nand2_1 U15419 ( .ip1(\pipeline/PC_DX [9]), .ip2(n18021), .op(n14261) );
  inv_1 U15420 ( .ip(n15896), .op(n20507) );
  nor2_1 U15421 ( .ip1(n20507), .ip2(n14392), .op(n14259) );
  nand2_1 U15422 ( .ip1(n14466), .ip2(\pipeline/epc [9]), .op(n14257) );
  nand2_1 U15423 ( .ip1(n10364), .ip2(\pipeline/csr/mtvec [9]), .op(n14256) );
  nand2_1 U15424 ( .ip1(n14257), .ip2(n14256), .op(n14258) );
  not_ab_or_c_or_d U15425 ( .ip1(\pipeline/PC_IF [9]), .ip2(n14404), .ip3(
        n14259), .ip4(n14258), .op(n14260) );
  nand2_1 U15426 ( .ip1(n14264), .ip2(n14263), .op(n14291) );
  xnor2_1 U15427 ( .ip1(n14264), .ip2(n14263), .op(n14585) );
  inv_1 U15428 ( .ip(n14265), .op(n14268) );
  inv_1 U15429 ( .ip(n14266), .op(n14267) );
  nand2_1 U15430 ( .ip1(n14268), .ip2(n14267), .op(n19687) );
  nor2_1 U15431 ( .ip1(n14274), .ip2(n14271), .op(n14284) );
  inv_1 U15432 ( .ip(n14272), .op(n14273) );
  nand2_1 U15433 ( .ip1(n14274), .ip2(n14273), .op(n14282) );
  nand2_1 U15434 ( .ip1(n10364), .ip2(\pipeline/csr/mtvec [11]), .op(n14277)
         );
  nand2_1 U15435 ( .ip1(n14282), .ip2(n14281), .op(n14283) );
  nor2_1 U15436 ( .ip1(n14284), .ip2(n14283), .op(n14293) );
  nand2_1 U15437 ( .ip1(n14285), .ip2(n14290), .op(n14294) );
  nand2_2 U15438 ( .ip1(n14288), .ip2(n14287), .op(n14308) );
  xor2_1 U15439 ( .ip1(n15308), .ip2(n14290), .op(n14292) );
  inv_1 U15440 ( .ip(n14293), .op(n14296) );
  inv_1 U15441 ( .ip(n14294), .op(n14295) );
  nand2_1 U15442 ( .ip1(n14296), .ip2(n14295), .op(n20689) );
  inv_1 U15443 ( .ip(n14300), .op(n14301) );
  nor2_1 U15444 ( .ip1(n14303), .ip2(n14225), .op(n14577) );
  inv_1 U15445 ( .ip(n14577), .op(n14304) );
  nand2_2 U15446 ( .ip1(n14309), .ip2(n17433), .op(n18299) );
  inv_1 U15447 ( .ip(\pipeline/PC_DX [20]), .op(n14311) );
  or2_1 U15448 ( .ip1(n14311), .ip2(n14310), .op(n14317) );
  inv_1 U15449 ( .ip(n15356), .op(n20584) );
  nor2_1 U15450 ( .ip1(n20584), .ip2(n14392), .op(n14315) );
  nand2_1 U15451 ( .ip1(n14466), .ip2(\pipeline/epc [20]), .op(n14313) );
  nand2_1 U15452 ( .ip1(n10364), .ip2(\pipeline/csr/mtvec [20]), .op(n14312)
         );
  nand2_1 U15453 ( .ip1(n14313), .ip2(n14312), .op(n14314) );
  not_ab_or_c_or_d U15454 ( .ip1(\pipeline/PC_IF [20]), .ip2(n14404), .ip3(
        n14315), .ip4(n14314), .op(n14316) );
  nand2_1 U15455 ( .ip1(n14317), .ip2(n14316), .op(n14379) );
  inv_1 U15456 ( .ip(n14379), .op(n14319) );
  and2_1 U15457 ( .ip1(n14318), .ip2(\pipeline/imm[31] ), .op(n14329) );
  inv_1 U15458 ( .ip(n14377), .op(n14320) );
  nand2_1 U15459 ( .ip1(\pipeline/PC_IF [19]), .ip2(n14404), .op(n14326) );
  nand2_1 U15460 ( .ip1(n14466), .ip2(\pipeline/epc [19]), .op(n14322) );
  nand2_1 U15461 ( .ip1(n10364), .ip2(\pipeline/csr/mtvec [19]), .op(n14321)
         );
  nand2_1 U15462 ( .ip1(n14322), .ip2(n14321), .op(n14324) );
  inv_1 U15463 ( .ip(n15628), .op(n20571) );
  nor2_1 U15464 ( .ip1(n20571), .ip2(n14392), .op(n14323) );
  nor2_1 U15465 ( .ip1(n14324), .ip2(n14323), .op(n14325) );
  nand2_1 U15466 ( .ip1(n14332), .ip2(n14327), .op(n14334) );
  nand2_1 U15467 ( .ip1(n14031), .ip2(\pipeline/inst_DX [19]), .op(n14328) );
  nand2_1 U15468 ( .ip1(n14334), .ip2(n14331), .op(n14381) );
  inv_1 U15469 ( .ip(n14329), .op(n14378) );
  nand2_1 U15470 ( .ip1(n14379), .ip2(n14378), .op(n14330) );
  inv_1 U15471 ( .ip(n14331), .op(n14333) );
  nand2_1 U15472 ( .ip1(n14031), .ip2(\pipeline/inst_DX [18]), .op(n14338) );
  inv_1 U15473 ( .ip(n15597), .op(n14609) );
  nor2_1 U15474 ( .ip1(n14609), .ip2(n14392), .op(n14344) );
  nand2_1 U15475 ( .ip1(n14466), .ip2(\pipeline/epc [18]), .op(n14342) );
  nand2_1 U15476 ( .ip1(n10364), .ip2(\pipeline/csr/mtvec [18]), .op(n14341)
         );
  nand2_1 U15477 ( .ip1(n14342), .ip2(n14341), .op(n14343) );
  nand2_1 U15478 ( .ip1(n14351), .ip2(n14350), .op(n14353) );
  nand2_1 U15479 ( .ip1(n14349), .ip2(n14348), .op(n14357) );
  inv_1 U15480 ( .ip(n14352), .op(n14355) );
  inv_1 U15481 ( .ip(n14353), .op(n14354) );
  nand2_2 U15482 ( .ip1(n14356), .ip2(n18294), .op(n19490) );
  nand2_1 U15483 ( .ip1(n14358), .ip2(n14357), .op(n20019) );
  nand2_1 U15484 ( .ip1(n18295), .ip2(n20019), .op(n14437) );
  inv_1 U15485 ( .ip(n14437), .op(n20041) );
  nor2_1 U15486 ( .ip1(n19490), .ip2(n20041), .op(n14359) );
  nand2_2 U15487 ( .ip1(n14360), .ip2(n10234), .op(n14509) );
  nor2_1 U15488 ( .ip1(n14362), .ip2(n14361), .op(n14518) );
  inv_1 U15489 ( .ip(n14518), .op(n18296) );
  nor2_1 U15490 ( .ip1(n19490), .ip2(n14518), .op(n14375) );
  nor2_2 U15491 ( .ip1(n14364), .ip2(n14363), .op(n19894) );
  inv_1 U15492 ( .ip(n14366), .op(n14369) );
  inv_1 U15493 ( .ip(n14367), .op(n14368) );
  nand2_1 U15494 ( .ip1(n14369), .ip2(n14368), .op(n19893) );
  nand2_1 U15495 ( .ip1(n14370), .ip2(n19893), .op(n14519) );
  nand2_1 U15496 ( .ip1(n14519), .ip2(n18285), .op(n14443) );
  inv_1 U15497 ( .ip(n14371), .op(n14372) );
  nor2_1 U15498 ( .ip1(n14373), .ip2(n14372), .op(n18287) );
  inv_1 U15499 ( .ip(n18287), .op(n14522) );
  nand2_1 U15500 ( .ip1(n14443), .ip2(n14522), .op(n14374) );
  nand2_1 U15501 ( .ip1(n14374), .ip2(n14440), .op(n18297) );
  nand2_1 U15502 ( .ip1(n14375), .ip2(n18297), .op(n14376) );
  nand2_1 U15503 ( .ip1(n14376), .ip2(n10234), .op(n14510) );
  inv_1 U15504 ( .ip(n14511), .op(n14386) );
  nand2_1 U15505 ( .ip1(n14377), .ip2(n14386), .op(n20036) );
  xnor2_1 U15506 ( .ip1(n14329), .ip2(n14379), .op(n14380) );
  inv_1 U15507 ( .ip(n14380), .op(n14383) );
  inv_1 U15508 ( .ip(n14381), .op(n14382) );
  nand2_1 U15509 ( .ip1(n14383), .ip2(n14382), .op(n19489) );
  nand2_2 U15510 ( .ip1(n14509), .ip2(n10215), .op(n14505) );
  nand2_1 U15511 ( .ip1(n14436), .ip2(n14505), .op(n14388) );
  inv_1 U15512 ( .ip(n14504), .op(n14506) );
  nand2_1 U15513 ( .ip1(n14386), .ip2(n14506), .op(n14451) );
  nand2_1 U15514 ( .ip1(n14451), .ip2(n14503), .op(n14387) );
  nand2_1 U15515 ( .ip1(n14388), .ip2(n14387), .op(n14389) );
  xor2_1 U15516 ( .ip1(n14511), .ip2(n14506), .op(n14391) );
  xor2_1 U15517 ( .ip1(n14391), .ip2(n14505), .op(imem_haddr[22]) );
  inv_1 U15518 ( .ip(n20650), .op(n21622) );
  nor2_1 U15519 ( .ip1(n21622), .ip2(n14392), .op(n14396) );
  nand2_1 U15520 ( .ip1(n14466), .ip2(\pipeline/epc [29]), .op(n14394) );
  nand2_1 U15521 ( .ip1(n10364), .ip2(\pipeline/csr/mtvec [29]), .op(n14393)
         );
  nand2_1 U15522 ( .ip1(n14394), .ip2(n14393), .op(n14395) );
  not_ab_or_c_or_d U15523 ( .ip1(\pipeline/PC_IF [29]), .ip2(n18024), .ip3(
        n14396), .ip4(n14395), .op(n14398) );
  nand2_1 U15524 ( .ip1(n14340), .ip2(\pipeline/PC_DX [29]), .op(n14397) );
  nand2_1 U15525 ( .ip1(n14398), .ip2(n14397), .op(n14546) );
  inv_1 U15526 ( .ip(n14546), .op(n14427) );
  nand2_1 U15527 ( .ip1(n14399), .ip2(\pipeline/PC_DX [25]), .op(n14406) );
  inv_1 U15528 ( .ip(n15565), .op(n20158) );
  nor2_1 U15529 ( .ip1(n20158), .ip2(n14392), .op(n14403) );
  nand2_1 U15530 ( .ip1(n14466), .ip2(\pipeline/epc [25]), .op(n14401) );
  nand2_1 U15531 ( .ip1(n10364), .ip2(\pipeline/csr/mtvec [25]), .op(n14400)
         );
  nand2_1 U15532 ( .ip1(n14401), .ip2(n14400), .op(n14402) );
  not_ab_or_c_or_d U15533 ( .ip1(\pipeline/PC_IF [25]), .ip2(n14404), .ip3(
        n14403), .ip4(n14402), .op(n14405) );
  nand2_1 U15534 ( .ip1(n14406), .ip2(n14405), .op(n14494) );
  nor2_1 U15535 ( .ip1(n14497), .ip2(n14494), .op(n14570) );
  nand2_1 U15536 ( .ip1(\pipeline/PC_DX [26]), .ip2(n14413), .op(n14412) );
  inv_1 U15537 ( .ip(n16333), .op(n16334) );
  nor2_1 U15538 ( .ip1(n16334), .ip2(n14392), .op(n14410) );
  nand2_1 U15539 ( .ip1(n14466), .ip2(\pipeline/epc [26]), .op(n14408) );
  nand2_1 U15540 ( .ip1(n10364), .ip2(\pipeline/csr/mtvec [26]), .op(n14407)
         );
  nand2_1 U15541 ( .ip1(n14408), .ip2(n14407), .op(n14409) );
  not_ab_or_c_or_d U15542 ( .ip1(\pipeline/PC_IF [26]), .ip2(n18024), .ip3(
        n14410), .ip4(n14409), .op(n14411) );
  and2_1 U15543 ( .ip1(n14412), .ip2(n14411), .op(n14568) );
  and2_1 U15544 ( .ip1(n14570), .ip2(n14568), .op(n14531) );
  nand2_1 U15545 ( .ip1(n14413), .ip2(\pipeline/PC_DX [27]), .op(n14419) );
  inv_1 U15546 ( .ip(n16237), .op(n16238) );
  nor2_1 U15547 ( .ip1(n16238), .ip2(n14392), .op(n14417) );
  nand2_1 U15548 ( .ip1(n14466), .ip2(\pipeline/epc [27]), .op(n14415) );
  nand2_1 U15549 ( .ip1(n10364), .ip2(\pipeline/csr/mtvec [27]), .op(n14414)
         );
  nand2_1 U15550 ( .ip1(n14415), .ip2(n14414), .op(n14416) );
  not_ab_or_c_or_d U15551 ( .ip1(\pipeline/PC_IF [27]), .ip2(n18024), .ip3(
        n14417), .ip4(n14416), .op(n14418) );
  nand2_1 U15552 ( .ip1(n14419), .ip2(n14418), .op(n14551) );
  nand2_1 U15553 ( .ip1(n14399), .ip2(\pipeline/PC_DX [28]), .op(n14425) );
  inv_1 U15554 ( .ip(n20646), .op(n20635) );
  nor2_1 U15555 ( .ip1(n20635), .ip2(n14392), .op(n14423) );
  nand2_1 U15556 ( .ip1(n14466), .ip2(\pipeline/epc [28]), .op(n14421) );
  nand2_1 U15557 ( .ip1(n10364), .ip2(\pipeline/csr/mtvec [28]), .op(n14420)
         );
  nand2_1 U15558 ( .ip1(n14421), .ip2(n14420), .op(n14422) );
  not_ab_or_c_or_d U15559 ( .ip1(\pipeline/PC_IF [28]), .ip2(n18024), .ip3(
        n14423), .ip4(n14422), .op(n14424) );
  nand2_1 U15560 ( .ip1(n14425), .ip2(n14424), .op(n14556) );
  nor2_1 U15561 ( .ip1(n14551), .ip2(n14556), .op(n14426) );
  nand2_1 U15562 ( .ip1(n14531), .ip2(n14426), .op(n14428) );
  nand2_1 U15563 ( .ip1(n14428), .ip2(n14427), .op(n14527) );
  inv_1 U15564 ( .ip(n14527), .op(n14429) );
  nor2_1 U15565 ( .ip1(n14546), .ip2(n14429), .op(n14459) );
  mux2_1 U15566 ( .ip1(n14568), .ip2(n14497), .s(n14494), .op(n14558) );
  nand2_1 U15567 ( .ip1(n14551), .ip2(n14556), .op(n14430) );
  nand2_1 U15568 ( .ip1(n14430), .ip2(n14546), .op(n14432) );
  nand2_1 U15569 ( .ip1(n14568), .ip2(n14551), .op(n14431) );
  and2_1 U15570 ( .ip1(n14432), .ip2(n14431), .op(n14433) );
  nand2_1 U15571 ( .ip1(n14558), .ip2(n14433), .op(n14434) );
  inv_1 U15572 ( .ip(n14434), .op(n14480) );
  nor2_1 U15573 ( .ip1(n14518), .ip2(n18287), .op(n14444) );
  inv_1 U15574 ( .ip(n14440), .op(n14517) );
  not_ab_or_c_or_d U15575 ( .ip1(n14444), .ip2(n14443), .ip3(n14442), .ip4(
        n14441), .op(n14456) );
  inv_1 U15576 ( .ip(n14448), .op(n14449) );
  nand2_1 U15577 ( .ip1(n14450), .ip2(n14449), .op(n14454) );
  inv_1 U15578 ( .ip(n14503), .op(n14452) );
  nor2_1 U15579 ( .ip1(n14452), .ip2(n14451), .op(n14453) );
  nand2_2 U15580 ( .ip1(n14458), .ip2(n14457), .op(n14532) );
  nand2_2 U15581 ( .ip1(n14480), .ip2(n14532), .op(n14528) );
  inv_1 U15582 ( .ip(n21645), .op(n21625) );
  nor2_1 U15583 ( .ip1(n21625), .ip2(n14392), .op(n14463) );
  nand2_1 U15584 ( .ip1(n14466), .ip2(\pipeline/epc [30]), .op(n14461) );
  nand2_1 U15585 ( .ip1(n10364), .ip2(\pipeline/csr/mtvec [30]), .op(n14460)
         );
  nand2_1 U15586 ( .ip1(n14461), .ip2(n14460), .op(n14462) );
  not_ab_or_c_or_d U15587 ( .ip1(\pipeline/PC_IF [30]), .ip2(n18024), .ip3(
        n14463), .ip4(n14462), .op(n14465) );
  nand2_1 U15588 ( .ip1(n18021), .ip2(\pipeline/PC_DX [30]), .op(n14464) );
  nand2_1 U15589 ( .ip1(n14465), .ip2(n14464), .op(n14526) );
  nand2_1 U15590 ( .ip1(n18021), .ip2(\pipeline/PC_DX [31]), .op(n14472) );
  inv_1 U15591 ( .ip(n14594), .op(n16020) );
  nor2_1 U15592 ( .ip1(n16020), .ip2(n14392), .op(n14470) );
  nand2_1 U15593 ( .ip1(n14466), .ip2(\pipeline/epc [31]), .op(n14468) );
  nand2_1 U15594 ( .ip1(n10364), .ip2(\pipeline/csr/mtvec [31]), .op(n14467)
         );
  nand2_1 U15595 ( .ip1(n14468), .ip2(n14467), .op(n14469) );
  not_ab_or_c_or_d U15596 ( .ip1(\pipeline/PC_IF [31]), .ip2(n18024), .ip3(
        n14470), .ip4(n14469), .op(n14471) );
  nand2_1 U15597 ( .ip1(n14472), .ip2(n14471), .op(n14473) );
  xor2_1 U15598 ( .ip1(n14473), .ip2(n14526), .op(n14483) );
  nor2_1 U15599 ( .ip1(n14526), .ip2(n14483), .op(n14474) );
  inv_1 U15600 ( .ip(n14483), .op(n14478) );
  inv_1 U15601 ( .ip(n14526), .op(n14479) );
  or2_1 U15602 ( .ip1(n14479), .ip2(n14478), .op(n14485) );
  nand2_1 U15603 ( .ip1(n14527), .ip2(n14483), .op(n14484) );
  nor2_1 U15604 ( .ip1(n14546), .ip2(n14484), .op(n14487) );
  inv_1 U15605 ( .ip(n14494), .op(n14498) );
  xor2_1 U15606 ( .ip1(n14497), .ip2(n14498), .op(n14493) );
  xor2_1 U15607 ( .ip1(n14494), .ip2(n14568), .op(n14502) );
  inv_1 U15608 ( .ip(n14497), .op(n14495) );
  nand2_1 U15609 ( .ip1(n14495), .ip2(n14494), .op(n14496) );
  nand2_1 U15610 ( .ip1(n14498), .ip2(n14497), .op(n14499) );
  nand2_2 U15611 ( .ip1(n14500), .ip2(n14499), .op(n14501) );
  xor2_2 U15612 ( .ip1(n14502), .ip2(n14501), .op(imem_haddr[26]) );
  xor2_1 U15613 ( .ip1(n14504), .ip2(n14503), .op(n14516) );
  nand3_1 U15614 ( .ip1(n14510), .ip2(n14509), .ip3(n14508), .op(n14512) );
  xor2_2 U15615 ( .ip1(n14516), .ip2(n14515), .op(imem_haddr[23]) );
  nor2_1 U15616 ( .ip1(n14518), .ip2(n14517), .op(n14525) );
  inv_1 U15617 ( .ip(n14519), .op(n14520) );
  xor2_2 U15618 ( .ip1(n14525), .ip2(n14524), .op(imem_haddr[17]) );
  xnor2_1 U15619 ( .ip1(n14526), .ip2(n14546), .op(n14530) );
  xor2_2 U15620 ( .ip1(n14530), .ip2(n14529), .op(imem_haddr[30]) );
  xor2_1 U15621 ( .ip1(n14551), .ip2(n14556), .op(n14539) );
  inv_1 U15622 ( .ip(n14539), .op(n14537) );
  inv_1 U15623 ( .ip(n14551), .op(n14567) );
  or2_1 U15624 ( .ip1(n14531), .ip2(n14551), .op(n14540) );
  nand2_1 U15625 ( .ip1(n14537), .ip2(n14540), .op(n14533) );
  nand2_2 U15626 ( .ip1(n14558), .ip2(n14532), .op(n14573) );
  or2_1 U15627 ( .ip1(n14533), .ip2(n14536), .op(n14545) );
  inv_1 U15628 ( .ip(n14568), .op(n14571) );
  nor2_1 U15629 ( .ip1(n14537), .ip2(n14534), .op(n14535) );
  nand2_1 U15630 ( .ip1(n14534), .ip2(n14537), .op(n14538) );
  nand2_1 U15631 ( .ip1(n14538), .ip2(n14540), .op(n14542) );
  or2_1 U15632 ( .ip1(n14540), .ip2(n14539), .op(n14541) );
  nand2_1 U15633 ( .ip1(n14542), .ip2(n14541), .op(n14543) );
  xor2_1 U15634 ( .ip1(n14546), .ip2(n14556), .op(n14559) );
  inv_1 U15635 ( .ip(n14559), .op(n14547) );
  nand2_1 U15636 ( .ip1(n14573), .ip2(n14548), .op(n14550) );
  nand2_1 U15637 ( .ip1(n14559), .ip2(n14556), .op(n14549) );
  nor2_1 U15638 ( .ip1(n14559), .ip2(n14556), .op(n14560) );
  and2_2 U15639 ( .ip1(n14566), .ip2(n10221), .op(imem_haddr[29]) );
  or2_1 U15640 ( .ip1(n14571), .ip2(n14570), .op(n14572) );
  xor2_2 U15641 ( .ip1(n14569), .ip2(n14574), .op(imem_haddr[27]) );
  nor2_1 U15642 ( .ip1(n14577), .ip2(n14576), .op(n14592) );
  inv_1 U15643 ( .ip(n14579), .op(n18309) );
  inv_1 U15644 ( .ip(n19688), .op(n14584) );
  inv_1 U15645 ( .ip(n14580), .op(n14581) );
  nand2_2 U15646 ( .ip1(n19689), .ip2(n19687), .op(n14583) );
  nand2_2 U15647 ( .ip1(n14584), .ip2(n14583), .op(n19763) );
  inv_1 U15648 ( .ip(n14585), .op(n19764) );
  nand2_2 U15649 ( .ip1(n19763), .ip2(n19764), .op(n18310) );
  nor2_2 U15650 ( .ip1(n18309), .ip2(n18310), .op(n20691) );
  nand2_1 U15651 ( .ip1(n20690), .ip2(n20691), .op(n14588) );
  inv_1 U15652 ( .ip(n14586), .op(n14587) );
  xor2_2 U15653 ( .ip1(n14592), .ip2(n14591), .op(imem_haddr[13]) );
  nor2_1 U15654 ( .ip1(n16478), .ip2(n15312), .op(n14595) );
  nor2_1 U15655 ( .ip1(n14596), .ip2(n14595), .op(n21646) );
  nand2_1 U15656 ( .ip1(n14594), .ip2(n21646), .op(n20483) );
  nor2_1 U15657 ( .ip1(n15467), .ip2(n20483), .op(n14606) );
  nor2_1 U15658 ( .ip1(n15433), .ip2(n20483), .op(n14600) );
  nor2_1 U15659 ( .ip1(n18022), .ip2(n14597), .op(n17344) );
  nand2_1 U15660 ( .ip1(n17344), .ip2(n17345), .op(n17853) );
  nor2_1 U15661 ( .ip1(n15796), .ip2(n17853), .op(n17938) );
  nand2_1 U15662 ( .ip1(n17938), .ip2(n15661), .op(n20474) );
  nor2_1 U15663 ( .ip1(n20476), .ip2(n20474), .op(n20484) );
  nand2_1 U15664 ( .ip1(n20484), .ip2(n15962), .op(n14598) );
  inv_1 U15665 ( .ip(n20483), .op(n21624) );
  nand2_1 U15666 ( .ip1(n14598), .ip2(n21624), .op(n20380) );
  nand2_1 U15667 ( .ip1(n21624), .ip2(n15928), .op(n14599) );
  nand2_1 U15668 ( .ip1(n20380), .ip2(n14599), .op(n19747) );
  nor2_1 U15669 ( .ip1(n14600), .ip2(n19747), .op(n20506) );
  nor2_1 U15670 ( .ip1(n20507), .ip2(n20483), .op(n14602) );
  nor2_1 U15671 ( .ip1(n14601), .ip2(n14602), .op(n14603) );
  and2_1 U15672 ( .ip1(n20506), .ip2(n14603), .op(n20522) );
  inv_1 U15673 ( .ip(n16226), .op(n20523) );
  nand2_1 U15674 ( .ip1(n20522), .ip2(n20523), .op(n14604) );
  nand2_1 U15675 ( .ip1(n14604), .ip2(n21624), .op(n20391) );
  nand2_1 U15676 ( .ip1(n21624), .ip2(n16402), .op(n14605) );
  nand2_1 U15677 ( .ip1(n20391), .ip2(n14605), .op(n20399) );
  nor2_1 U15678 ( .ip1(n14606), .ip2(n20399), .op(n20423) );
  nor2_1 U15679 ( .ip1(n20424), .ip2(n20483), .op(n14607) );
  nor2_1 U15680 ( .ip1(n20426), .ip2(n14607), .op(n14608) );
  nand2_1 U15681 ( .ip1(n20423), .ip2(n14608), .op(n20430) );
  nor2_1 U15682 ( .ip1(n14593), .ip2(n20430), .op(n20005) );
  and2_1 U15683 ( .ip1(n20005), .ip2(n15499), .op(n20440) );
  nand2_1 U15684 ( .ip1(n20440), .ip2(n14609), .op(n14610) );
  nand2_1 U15685 ( .ip1(n14610), .ip2(n21624), .op(n20570) );
  nand2_1 U15686 ( .ip1(n20570), .ip2(n20571), .op(n14611) );
  nand2_1 U15687 ( .ip1(n14611), .ip2(n21624), .op(n20583) );
  nor2_1 U15688 ( .ip1(n20584), .ip2(n20483), .op(n14612) );
  nor2_1 U15689 ( .ip1(n20586), .ip2(n14612), .op(n14613) );
  nand2_1 U15690 ( .ip1(n20583), .ip2(n14613), .op(n20598) );
  nor2_1 U15691 ( .ip1(n15369), .ip2(n20598), .op(n20277) );
  and2_1 U15692 ( .ip1(n20277), .ip2(n20278), .op(n20609) );
  nand2_1 U15693 ( .ip1(n20609), .ip2(n16112), .op(n14614) );
  nand2_1 U15694 ( .ip1(n14614), .ip2(n21624), .op(n20157) );
  and2_1 U15695 ( .ip1(n20157), .ip2(n20158), .op(n20622) );
  nand2_1 U15696 ( .ip1(n20622), .ip2(n16334), .op(n14772) );
  nand2_1 U15697 ( .ip1(n14772), .ip2(n21624), .op(n14615) );
  nand2_1 U15698 ( .ip1(n14615), .ip2(n16238), .op(n20645) );
  or2_1 U15699 ( .ip1(n17788), .ip2(n17819), .op(n21683) );
  inv_1 U15700 ( .ip(\pipeline/md/a [46]), .op(n21851) );
  nor2_1 U15701 ( .ip1(\pipeline/md/b [46]), .ip2(n21851), .op(n14616) );
  inv_1 U15702 ( .ip(\pipeline/md/a [45]), .op(n14721) );
  nor2_1 U15703 ( .ip1(\pipeline/md/b [45]), .ip2(n14721), .op(n21846) );
  nor2_1 U15704 ( .ip1(n14616), .ip2(n21846), .op(n21708) );
  inv_1 U15705 ( .ip(\pipeline/md/b [44]), .op(n14617) );
  nand2_1 U15706 ( .ip1(\pipeline/md/a [44]), .ip2(n14617), .op(n21832) );
  inv_1 U15707 ( .ip(\pipeline/md/a [43]), .op(n14618) );
  nor2_1 U15708 ( .ip1(\pipeline/md/b [43]), .ip2(n14618), .op(n21824) );
  inv_1 U15709 ( .ip(\pipeline/md/b [42]), .op(n21822) );
  nor2_1 U15710 ( .ip1(\pipeline/md/a [42]), .ip2(n21822), .op(n14619) );
  inv_1 U15711 ( .ip(\pipeline/md/b [43]), .op(n21390) );
  nor2_1 U15712 ( .ip1(\pipeline/md/a [43]), .ip2(n21390), .op(n21823) );
  nor2_1 U15713 ( .ip1(n14619), .ip2(n21823), .op(n14620) );
  nor2_1 U15714 ( .ip1(n21824), .ip2(n14620), .op(n14628) );
  inv_1 U15715 ( .ip(\pipeline/md/b [40]), .op(n21758) );
  nor2_1 U15716 ( .ip1(\pipeline/md/a [40]), .ip2(n21758), .op(n14622) );
  inv_1 U15717 ( .ip(\pipeline/md/b [41]), .op(n21763) );
  nor2_1 U15718 ( .ip1(\pipeline/md/a [41]), .ip2(n21763), .op(n14621) );
  nor2_1 U15719 ( .ip1(n14622), .ip2(n14621), .op(n14626) );
  inv_1 U15720 ( .ip(n21824), .op(n14625) );
  nand2_1 U15721 ( .ip1(\pipeline/md/a [42]), .ip2(n21822), .op(n14624) );
  nand2_1 U15722 ( .ip1(\pipeline/md/a [41]), .ip2(n21763), .op(n14623) );
  nand3_1 U15723 ( .ip1(n14625), .ip2(n14624), .ip3(n14623), .op(n21703) );
  nor2_1 U15724 ( .ip1(n14626), .ip2(n21703), .op(n14627) );
  or2_1 U15725 ( .ip1(n14628), .ip2(n14627), .op(n21705) );
  nand2_1 U15726 ( .ip1(n21832), .ip2(n21705), .op(n14723) );
  inv_1 U15727 ( .ip(n21703), .op(n14720) );
  inv_1 U15728 ( .ip(\pipeline/md/a [39]), .op(n14629) );
  nand2_1 U15729 ( .ip1(\pipeline/md/b [39]), .ip2(n14629), .op(n21692) );
  nor2_1 U15730 ( .ip1(\pipeline/md/b [39]), .ip2(n14629), .op(n21812) );
  inv_1 U15731 ( .ip(\pipeline/md/a [38]), .op(n14713) );
  nor2_1 U15732 ( .ip1(\pipeline/md/b [38]), .ip2(n14713), .op(n21805) );
  nor2_1 U15733 ( .ip1(n21812), .ip2(n21805), .op(n21701) );
  inv_1 U15734 ( .ip(\pipeline/md/a [35]), .op(n21783) );
  nor2_1 U15735 ( .ip1(\pipeline/md/b [35]), .ip2(n21783), .op(n14711) );
  inv_1 U15736 ( .ip(\pipeline/md/a [34]), .op(n21773) );
  inv_1 U15737 ( .ip(\pipeline/md/b [33]), .op(n22495) );
  nand2_1 U15738 ( .ip1(\pipeline/md/a [33]), .ip2(n22495), .op(n21799) );
  inv_1 U15739 ( .ip(\pipeline/md/a [32]), .op(n21791) );
  nand2_1 U15740 ( .ip1(\pipeline/md/b [32]), .ip2(n21791), .op(n21797) );
  or2_1 U15741 ( .ip1(\pipeline/md/a [33]), .ip2(n22495), .op(n21798) );
  nand2_1 U15742 ( .ip1(n21797), .ip2(n21798), .op(n14630) );
  and2_1 U15743 ( .ip1(n21799), .ip2(n14630), .op(n21693) );
  inv_1 U15744 ( .ip(\pipeline/md/b [32]), .op(n22484) );
  nand2_1 U15745 ( .ip1(\pipeline/md/a [32]), .ip2(n22484), .op(n21794) );
  inv_1 U15746 ( .ip(n21794), .op(n14703) );
  inv_1 U15747 ( .ip(n21799), .op(n14702) );
  inv_1 U15748 ( .ip(\pipeline/md/a [30]), .op(n14890) );
  nor2_1 U15749 ( .ip1(\pipeline/md/b [30]), .ip2(n14890), .op(n21639) );
  inv_1 U15750 ( .ip(n21639), .op(n14632) );
  inv_1 U15751 ( .ip(\pipeline/md/b [31]), .op(n21656) );
  nand2_1 U15752 ( .ip1(\pipeline/md/a [31]), .ip2(n21656), .op(n14631) );
  nand2_1 U15753 ( .ip1(n14632), .ip2(n14631), .op(n21694) );
  inv_1 U15754 ( .ip(n21694), .op(n14633) );
  nor2_1 U15755 ( .ip1(\pipeline/md/a [31]), .ip2(n21656), .op(n21697) );
  or2_1 U15756 ( .ip1(n14633), .ip2(n21697), .op(n14700) );
  inv_1 U15757 ( .ip(\pipeline/md/b [29]), .op(n20657) );
  nand2_1 U15758 ( .ip1(\pipeline/md/a [29]), .ip2(n20657), .op(n21630) );
  inv_1 U15759 ( .ip(\pipeline/md/b [28]), .op(n18844) );
  nor2_1 U15760 ( .ip1(\pipeline/md/a [28]), .ip2(n18844), .op(n20655) );
  inv_1 U15761 ( .ip(\pipeline/md/a [28]), .op(n14634) );
  nor2_1 U15762 ( .ip1(\pipeline/md/b [28]), .ip2(n14634), .op(n20653) );
  inv_1 U15763 ( .ip(\pipeline/md/b [26]), .op(n15273) );
  nand2_1 U15764 ( .ip1(\pipeline/md/a [26]), .ip2(n15273), .op(n14802) );
  inv_1 U15765 ( .ip(n14802), .op(n14691) );
  inv_1 U15766 ( .ip(\pipeline/md/a [27]), .op(n14822) );
  nor2_1 U15767 ( .ip1(\pipeline/md/b [27]), .ip2(n14822), .op(n14808) );
  inv_1 U15768 ( .ip(\pipeline/md/b [25]), .op(n15249) );
  nand2_1 U15769 ( .ip1(\pipeline/md/a [25]), .ip2(n15249), .op(n20150) );
  inv_1 U15770 ( .ip(\pipeline/md/a [24]), .op(n20617) );
  nand2_1 U15771 ( .ip1(\pipeline/md/b [24]), .ip2(n20617), .op(n14800) );
  inv_1 U15772 ( .ip(\pipeline/md/b [24]), .op(n20615) );
  nand2_1 U15773 ( .ip1(\pipeline/md/a [24]), .ip2(n20615), .op(n14797) );
  inv_1 U15774 ( .ip(\pipeline/md/b [22]), .op(n20602) );
  nor2_1 U15775 ( .ip1(\pipeline/md/a [22]), .ip2(n20602), .op(n20283) );
  inv_1 U15776 ( .ip(\pipeline/md/b [23]), .op(n15242) );
  nor2_1 U15777 ( .ip1(\pipeline/md/a [23]), .ip2(n15242), .op(n14635) );
  nor2_1 U15778 ( .ip1(n20283), .ip2(n14635), .op(n14637) );
  inv_1 U15779 ( .ip(\pipeline/md/a [23]), .op(n14636) );
  nor2_1 U15780 ( .ip1(\pipeline/md/b [23]), .ip2(n14636), .op(n14681) );
  nor2_1 U15781 ( .ip1(n14637), .ip2(n14681), .op(n14795) );
  inv_1 U15782 ( .ip(\pipeline/md/a [20]), .op(n14885) );
  nor2_1 U15783 ( .ip1(\pipeline/md/b [20]), .ip2(n14885), .op(n14792) );
  inv_1 U15784 ( .ip(n14792), .op(n14679) );
  inv_1 U15785 ( .ip(\pipeline/md/b [20]), .op(n20577) );
  nor2_1 U15786 ( .ip1(\pipeline/md/a [20]), .ip2(n20577), .op(n14790) );
  inv_1 U15787 ( .ip(n14790), .op(n14646) );
  inv_1 U15788 ( .ip(\pipeline/md/a [19]), .op(n14638) );
  nand2_1 U15789 ( .ip1(\pipeline/md/b [19]), .ip2(n14638), .op(n14788) );
  inv_1 U15790 ( .ip(\pipeline/md/b [18]), .op(n15194) );
  nand2_1 U15791 ( .ip1(\pipeline/md/a [18]), .ip2(n15194), .op(n20564) );
  inv_1 U15792 ( .ip(\pipeline/md/b [19]), .op(n15227) );
  nand2_1 U15793 ( .ip1(\pipeline/md/a [19]), .ip2(n15227), .op(n14642) );
  and2_1 U15794 ( .ip1(n20564), .ip2(n14642), .op(n14787) );
  inv_1 U15795 ( .ip(\pipeline/md/b [17]), .op(n20010) );
  nand2_1 U15796 ( .ip1(\pipeline/md/a [17]), .ip2(n20010), .op(n14785) );
  and2_1 U15797 ( .ip1(n14787), .ip2(n14785), .op(n14674) );
  inv_1 U15798 ( .ip(\pipeline/md/a [17]), .op(n14639) );
  nand2_1 U15799 ( .ip1(\pipeline/md/b [17]), .ip2(n14639), .op(n14783) );
  inv_1 U15800 ( .ip(\pipeline/md/b [16]), .op(n15166) );
  nor2_1 U15801 ( .ip1(\pipeline/md/a [16]), .ip2(n15166), .op(n14782) );
  inv_1 U15802 ( .ip(n14782), .op(n14640) );
  nand2_1 U15803 ( .ip1(n14783), .ip2(n14640), .op(n14641) );
  nand2_1 U15804 ( .ip1(n14674), .ip2(n14641), .op(n14645) );
  inv_1 U15805 ( .ip(\pipeline/md/a [18]), .op(n14824) );
  nand2_1 U15806 ( .ip1(\pipeline/md/b [18]), .ip2(n14824), .op(n14786) );
  inv_1 U15807 ( .ip(n14786), .op(n14643) );
  nand2_1 U15808 ( .ip1(n14643), .ip2(n14642), .op(n14644) );
  nand4_1 U15809 ( .ip1(n14646), .ip2(n14788), .ip3(n14645), .ip4(n14644), 
        .op(n14678) );
  inv_1 U15810 ( .ip(\pipeline/md/b [14]), .op(n20417) );
  nor2_1 U15811 ( .ip1(\pipeline/md/a [14]), .ip2(n20417), .op(n20433) );
  inv_1 U15812 ( .ip(\pipeline/md/b [15]), .op(n15144) );
  nor2_1 U15813 ( .ip1(\pipeline/md/a [15]), .ip2(n15144), .op(n14647) );
  nor2_1 U15814 ( .ip1(n20433), .ip2(n14647), .op(n14777) );
  inv_1 U15815 ( .ip(\pipeline/md/a [13]), .op(n14649) );
  nor2_1 U15816 ( .ip1(\pipeline/md/b [13]), .ip2(n14649), .op(n20411) );
  nand2_1 U15817 ( .ip1(\pipeline/md/b [13]), .ip2(n14649), .op(n20414) );
  inv_1 U15818 ( .ip(\pipeline/md/a [12]), .op(n14868) );
  nand2_1 U15819 ( .ip1(\pipeline/md/b [12]), .ip2(n14868), .op(n20402) );
  nand2_1 U15820 ( .ip1(n20414), .ip2(n20402), .op(n14671) );
  inv_1 U15821 ( .ip(\pipeline/md/b [10]), .op(n20515) );
  nor2_1 U15822 ( .ip1(\pipeline/md/a [10]), .ip2(n20515), .op(n20526) );
  inv_1 U15823 ( .ip(\pipeline/md/b [11]), .op(n15088) );
  nand2_1 U15824 ( .ip1(\pipeline/md/a [11]), .ip2(n15088), .op(n14669) );
  nor2_1 U15825 ( .ip1(\pipeline/md/a [11]), .ip2(n15088), .op(n14668) );
  inv_1 U15826 ( .ip(\pipeline/md/a [9]), .op(n14857) );
  nor2_1 U15827 ( .ip1(\pipeline/md/b [9]), .ip2(n14857), .op(n20514) );
  inv_1 U15828 ( .ip(\pipeline/md/b [8]), .op(n19756) );
  nand2_1 U15829 ( .ip1(\pipeline/md/a [8]), .ip2(n19756), .op(n20495) );
  inv_1 U15830 ( .ip(n20495), .op(n14661) );
  inv_1 U15831 ( .ip(\pipeline/md/a [6]), .op(n14873) );
  nand2_1 U15832 ( .ip1(\pipeline/md/b [6]), .ip2(n14873), .op(n19752) );
  inv_1 U15833 ( .ip(\pipeline/md/a [7]), .op(n14650) );
  nand2_1 U15834 ( .ip1(\pipeline/md/b [7]), .ip2(n14650), .op(n19755) );
  nand2_1 U15835 ( .ip1(n19752), .ip2(n19755), .op(n14659) );
  nor2_1 U15836 ( .ip1(\pipeline/md/b [6]), .ip2(n14873), .op(n14658) );
  inv_1 U15837 ( .ip(\pipeline/md/b [3]), .op(n17851) );
  inv_1 U15838 ( .ip(\pipeline/md/b [2]), .op(n17341) );
  inv_1 U15839 ( .ip(\pipeline/md/b [1]), .op(n17331) );
  inv_1 U15840 ( .ip(\pipeline/md/a [0]), .op(n14832) );
  nand2_1 U15841 ( .ip1(\pipeline/md/b [0]), .ip2(n14832), .op(n21501) );
  inv_1 U15842 ( .ip(\pipeline/md/b [4]), .op(n14936) );
  nor2_1 U15843 ( .ip1(n14651), .ip2(n14936), .op(n17943) );
  inv_1 U15844 ( .ip(n14651), .op(n14652) );
  nor2_1 U15845 ( .ip1(\pipeline/md/b [4]), .ip2(n14652), .op(n17942) );
  nor2_1 U15846 ( .ip1(\pipeline/md/a [4]), .ip2(n17942), .op(n14653) );
  nor2_1 U15847 ( .ip1(n17943), .ip2(n14653), .op(n20479) );
  inv_1 U15848 ( .ip(\pipeline/md/a [5]), .op(n14654) );
  nand2_1 U15849 ( .ip1(\pipeline/md/b [5]), .ip2(n14654), .op(n14655) );
  nand2_1 U15850 ( .ip1(n20479), .ip2(n14655), .op(n14657) );
  inv_1 U15851 ( .ip(\pipeline/md/b [5]), .op(n14965) );
  nand2_1 U15852 ( .ip1(\pipeline/md/a [5]), .ip2(n14965), .op(n14656) );
  nand2_1 U15853 ( .ip1(n14657), .ip2(n14656), .op(n20488) );
  nor2_1 U15854 ( .ip1(n14658), .ip2(n20488), .op(n19750) );
  nor2_1 U15855 ( .ip1(n14659), .ip2(n19750), .op(n14660) );
  nor2_1 U15856 ( .ip1(n14661), .ip2(n14660), .op(n14665) );
  inv_1 U15857 ( .ip(\pipeline/md/b [7]), .op(n14662) );
  nand2_1 U15858 ( .ip1(\pipeline/md/a [7]), .ip2(n14662), .op(n19753) );
  inv_1 U15859 ( .ip(\pipeline/md/b [9]), .op(n20500) );
  nor2_1 U15860 ( .ip1(\pipeline/md/a [9]), .ip2(n20500), .op(n14664) );
  inv_1 U15861 ( .ip(\pipeline/md/a [8]), .op(n14829) );
  nand2_1 U15862 ( .ip1(\pipeline/md/b [8]), .ip2(n14829), .op(n20497) );
  inv_1 U15863 ( .ip(n20497), .op(n14663) );
  not_ab_or_c_or_d U15864 ( .ip1(n14665), .ip2(n19753), .ip3(n14664), .ip4(
        n14663), .op(n20513) );
  nand2_1 U15865 ( .ip1(\pipeline/md/a [10]), .ip2(n20515), .op(n20528) );
  nand2_1 U15866 ( .ip1(n20528), .ip2(n14669), .op(n14666) );
  nor3_1 U15867 ( .ip1(n20514), .ip2(n20513), .ip3(n14666), .op(n14667) );
  not_ab_or_c_or_d U15868 ( .ip1(n20526), .ip2(n14669), .ip3(n14668), .ip4(
        n14667), .op(n20403) );
  nor2_1 U15869 ( .ip1(\pipeline/md/b [12]), .ip2(n14868), .op(n20412) );
  nor2_1 U15870 ( .ip1(n20403), .ip2(n20412), .op(n14670) );
  nor2_1 U15871 ( .ip1(n14671), .ip2(n14670), .op(n14672) );
  or3_1 U15872 ( .ip1(n14648), .ip2(n20411), .ip3(n14672), .op(n20431) );
  inv_1 U15873 ( .ip(\pipeline/md/a [15]), .op(n14673) );
  nor2_1 U15874 ( .ip1(\pipeline/md/b [15]), .ip2(n14673), .op(n14776) );
  inv_1 U15875 ( .ip(\pipeline/md/a [16]), .op(n14826) );
  nor2_1 U15876 ( .ip1(\pipeline/md/b [16]), .ip2(n14826), .op(n14780) );
  or3_1 U15877 ( .ip1(n14776), .ip2(n14792), .ip3(n14780), .op(n14676) );
  inv_1 U15878 ( .ip(n14674), .op(n14675) );
  not_ab_or_c_or_d U15879 ( .ip1(n14777), .ip2(n20431), .ip3(n14676), .ip4(
        n14675), .op(n14677) );
  inv_1 U15880 ( .ip(\pipeline/md/b [21]), .op(n20590) );
  nor2_1 U15881 ( .ip1(\pipeline/md/a [21]), .ip2(n20590), .op(n14793) );
  not_ab_or_c_or_d U15882 ( .ip1(n14679), .ip2(n14678), .ip3(n14677), .ip4(
        n14793), .op(n14682) );
  inv_1 U15883 ( .ip(\pipeline/md/a [22]), .op(n14886) );
  nor2_1 U15884 ( .ip1(\pipeline/md/b [22]), .ip2(n14886), .op(n20285) );
  inv_1 U15885 ( .ip(\pipeline/md/a [21]), .op(n14680) );
  nor2_1 U15886 ( .ip1(\pipeline/md/b [21]), .ip2(n14680), .op(n20281) );
  or3_1 U15887 ( .ip1(n14681), .ip2(n20285), .ip3(n20281), .op(n14794) );
  nor2_1 U15888 ( .ip1(n14682), .ip2(n14794), .op(n14683) );
  or2_1 U15889 ( .ip1(n14795), .ip2(n14683), .op(n14684) );
  nand2_1 U15890 ( .ip1(n14797), .ip2(n14684), .op(n14685) );
  nand2_1 U15891 ( .ip1(n14800), .ip2(n14685), .op(n14689) );
  inv_1 U15892 ( .ip(\pipeline/md/a [26]), .op(n14686) );
  nand2_1 U15893 ( .ip1(\pipeline/md/b [26]), .ip2(n14686), .op(n14804) );
  inv_1 U15894 ( .ip(n14804), .op(n14688) );
  nor2_1 U15895 ( .ip1(\pipeline/md/a [25]), .ip2(n15249), .op(n14687) );
  not_ab_or_c_or_d U15896 ( .ip1(n20150), .ip2(n14689), .ip3(n14688), .ip4(
        n14687), .op(n14690) );
  nor3_1 U15897 ( .ip1(n14691), .ip2(n14808), .ip3(n14690), .op(n14693) );
  inv_1 U15898 ( .ip(\pipeline/md/b [27]), .op(n15279) );
  nor2_1 U15899 ( .ip1(\pipeline/md/a [27]), .ip2(n15279), .op(n14692) );
  nor2_1 U15900 ( .ip1(n14693), .ip2(n14692), .op(n14694) );
  nor2_1 U15901 ( .ip1(n20653), .ip2(n14694), .op(n14695) );
  or2_1 U15902 ( .ip1(n20655), .ip2(n14695), .op(n14697) );
  inv_1 U15903 ( .ip(\pipeline/md/b [30]), .op(n18850) );
  nor2_1 U15904 ( .ip1(\pipeline/md/a [30]), .ip2(n18850), .op(n21637) );
  inv_1 U15905 ( .ip(\pipeline/md/a [29]), .op(n14820) );
  nand2_1 U15906 ( .ip1(\pipeline/md/b [29]), .ip2(n14820), .op(n21627) );
  inv_1 U15907 ( .ip(n21627), .op(n14696) );
  ab_or_c_or_d U15908 ( .ip1(n21630), .ip2(n14697), .ip3(n21637), .ip4(n14696), 
        .op(n14698) );
  or2_1 U15909 ( .ip1(n14698), .ip2(n21697), .op(n14699) );
  nand2_1 U15910 ( .ip1(n14700), .ip2(n14699), .op(n14701) );
  nor3_1 U15911 ( .ip1(n14703), .ip2(n14702), .ip3(n14701), .op(n14704) );
  nor2_1 U15912 ( .ip1(n21693), .ip2(n14704), .op(n14706) );
  nor2_1 U15913 ( .ip1(\pipeline/md/b [34]), .ip2(n21773), .op(n14705) );
  nor2_1 U15914 ( .ip1(n14706), .ip2(n14705), .op(n14708) );
  inv_1 U15915 ( .ip(\pipeline/md/b [35]), .op(n21425) );
  nor2_1 U15916 ( .ip1(\pipeline/md/a [35]), .ip2(n21425), .op(n14707) );
  not_ab_or_c_or_d U15917 ( .ip1(\pipeline/md/b [34]), .ip2(n21773), .ip3(
        n14708), .ip4(n14707), .op(n14710) );
  inv_1 U15918 ( .ip(\pipeline/md/a [36]), .op(n21768) );
  nor2_1 U15919 ( .ip1(\pipeline/md/b [36]), .ip2(n21768), .op(n14709) );
  inv_1 U15920 ( .ip(\pipeline/md/a [37]), .op(n21778) );
  nor2_1 U15921 ( .ip1(\pipeline/md/b [37]), .ip2(n21778), .op(n14712) );
  or4_1 U15922 ( .ip1(n14711), .ip2(n14710), .ip3(n14709), .ip4(n14712), .op(
        n14716) );
  inv_1 U15923 ( .ip(\pipeline/md/b [36]), .op(n17301) );
  or3_1 U15924 ( .ip1(n14712), .ip2(\pipeline/md/a [36]), .ip3(n17301), .op(
        n14715) );
  nand2_1 U15925 ( .ip1(\pipeline/md/b [38]), .ip2(n14713), .op(n21806) );
  nand2_1 U15926 ( .ip1(\pipeline/md/b [37]), .ip2(n21778), .op(n14714) );
  nand4_1 U15927 ( .ip1(n14716), .ip2(n14715), .ip3(n21806), .ip4(n14714), 
        .op(n14717) );
  nand2_1 U15928 ( .ip1(n21701), .ip2(n14717), .op(n14718) );
  nand2_1 U15929 ( .ip1(n21692), .ip2(n14718), .op(n14719) );
  nand2_1 U15930 ( .ip1(\pipeline/md/a [40]), .ip2(n21758), .op(n21691) );
  nand4_1 U15931 ( .ip1(n14720), .ip2(n21832), .ip3(n14719), .ip4(n21691), 
        .op(n14722) );
  inv_1 U15932 ( .ip(\pipeline/md/a [44]), .op(n21830) );
  nand2_1 U15933 ( .ip1(\pipeline/md/b [44]), .ip2(n21830), .op(n21831) );
  nand2_1 U15934 ( .ip1(\pipeline/md/b [45]), .ip2(n14721), .op(n21839) );
  nand4_1 U15935 ( .ip1(n14723), .ip2(n14722), .ip3(n21831), .ip4(n21839), 
        .op(n14725) );
  inv_1 U15936 ( .ip(\pipeline/md/b [47]), .op(n22619) );
  nor2_1 U15937 ( .ip1(\pipeline/md/a [47]), .ip2(n22619), .op(n21689) );
  inv_1 U15938 ( .ip(\pipeline/md/b [46]), .op(n14724) );
  nor2_1 U15939 ( .ip1(\pipeline/md/a [46]), .ip2(n14724), .op(n21690) );
  not_ab_or_c_or_d U15940 ( .ip1(n21708), .ip2(n14725), .ip3(n21689), .ip4(
        n21690), .op(n14729) );
  inv_1 U15941 ( .ip(\pipeline/md/b [53]), .op(n22680) );
  nand2_1 U15942 ( .ip1(\pipeline/md/a [53]), .ip2(n22680), .op(n21878) );
  inv_1 U15943 ( .ip(\pipeline/md/b [52]), .op(n14738) );
  nand2_1 U15944 ( .ip1(\pipeline/md/a [52]), .ip2(n14738), .op(n21874) );
  nand2_1 U15945 ( .ip1(n21878), .ip2(n21874), .op(n21717) );
  inv_1 U15946 ( .ip(\pipeline/md/b [54]), .op(n22690) );
  nand2_1 U15947 ( .ip1(\pipeline/md/a [54]), .ip2(n22690), .op(n21891) );
  inv_1 U15948 ( .ip(\pipeline/md/b [55]), .op(n22699) );
  nand2_1 U15949 ( .ip1(\pipeline/md/a [55]), .ip2(n22699), .op(n21896) );
  nand2_1 U15950 ( .ip1(n21891), .ip2(n21896), .op(n21720) );
  inv_1 U15951 ( .ip(\pipeline/md/b [50]), .op(n22650) );
  inv_1 U15952 ( .ip(\pipeline/md/a [51]), .op(n21745) );
  nor2_1 U15953 ( .ip1(\pipeline/md/b [51]), .ip2(n21745), .op(n14732) );
  inv_1 U15954 ( .ip(\pipeline/md/a [49]), .op(n21750) );
  nor2_1 U15955 ( .ip1(\pipeline/md/b [49]), .ip2(n21750), .op(n14726) );
  not_ab_or_c_or_d U15956 ( .ip1(\pipeline/md/a [50]), .ip2(n22650), .ip3(
        n14732), .ip4(n14726), .op(n14736) );
  inv_1 U15957 ( .ip(\pipeline/md/b [48]), .op(n22629) );
  nand2_1 U15958 ( .ip1(\pipeline/md/a [48]), .ip2(n22629), .op(n21714) );
  nand2_1 U15959 ( .ip1(\pipeline/md/a [47]), .ip2(n22619), .op(n21711) );
  inv_1 U15960 ( .ip(\pipeline/md/a [56]), .op(n21910) );
  nor2_1 U15961 ( .ip1(\pipeline/md/b [56]), .ip2(n21910), .op(n21904) );
  inv_1 U15962 ( .ip(\pipeline/md/a [57]), .op(n21922) );
  nor2_1 U15963 ( .ip1(\pipeline/md/b [57]), .ip2(n21922), .op(n21918) );
  or2_1 U15964 ( .ip1(n21904), .ip2(n21918), .op(n14746) );
  inv_1 U15965 ( .ip(n14746), .op(n14727) );
  nand4_1 U15966 ( .ip1(n14736), .ip2(n21714), .ip3(n21711), .ip4(n14727), 
        .op(n14728) );
  nor4_1 U15967 ( .ip1(n14729), .ip2(n21717), .ip3(n21720), .ip4(n14728), .op(
        n14748) );
  inv_1 U15968 ( .ip(n21720), .op(n14744) );
  inv_1 U15969 ( .ip(\pipeline/md/a [48]), .op(n14730) );
  nand2_1 U15970 ( .ip1(\pipeline/md/b [48]), .ip2(n14730), .op(n21716) );
  nand2_1 U15971 ( .ip1(\pipeline/md/b [49]), .ip2(n21750), .op(n14731) );
  nand2_1 U15972 ( .ip1(n21716), .ip2(n14731), .op(n14735) );
  inv_1 U15973 ( .ip(\pipeline/md/b [51]), .op(n21345) );
  nor2_1 U15974 ( .ip1(\pipeline/md/a [51]), .ip2(n21345), .op(n14734) );
  nor3_1 U15975 ( .ip1(n14732), .ip2(\pipeline/md/a [50]), .ip3(n22650), .op(
        n14733) );
  not_ab_or_c_or_d U15976 ( .ip1(n14736), .ip2(n14735), .ip3(n14734), .ip4(
        n14733), .op(n14737) );
  or2_1 U15977 ( .ip1(n14737), .ip2(n21717), .op(n14742) );
  nor2_1 U15978 ( .ip1(\pipeline/md/a [52]), .ip2(n14738), .op(n21867) );
  nand2_1 U15979 ( .ip1(n21867), .ip2(n21878), .op(n14741) );
  inv_1 U15980 ( .ip(\pipeline/md/a [54]), .op(n14739) );
  nand2_1 U15981 ( .ip1(\pipeline/md/b [54]), .ip2(n14739), .op(n21885) );
  inv_1 U15982 ( .ip(\pipeline/md/a [53]), .op(n14740) );
  nand2_1 U15983 ( .ip1(\pipeline/md/b [53]), .ip2(n14740), .op(n21877) );
  nand4_1 U15984 ( .ip1(n14742), .ip2(n14741), .ip3(n21885), .ip4(n21877), 
        .op(n14743) );
  inv_1 U15985 ( .ip(\pipeline/md/b [56]), .op(n21905) );
  nor2_1 U15986 ( .ip1(\pipeline/md/a [56]), .ip2(n21905), .op(n21723) );
  nor2_1 U15987 ( .ip1(\pipeline/md/a [55]), .ip2(n22699), .op(n21894) );
  not_ab_or_c_or_d U15988 ( .ip1(n14744), .ip2(n14743), .ip3(n21723), .ip4(
        n21894), .op(n14745) );
  nor2_1 U15989 ( .ip1(n14746), .ip2(n14745), .op(n14747) );
  inv_1 U15990 ( .ip(\pipeline/md/b [57]), .op(n21320) );
  nor2_1 U15991 ( .ip1(\pipeline/md/a [57]), .ip2(n21320), .op(n21725) );
  nor3_1 U15992 ( .ip1(n14748), .ip2(n14747), .ip3(n21725), .op(n14754) );
  inv_1 U15993 ( .ip(\pipeline/md/a [62]), .op(n21951) );
  nor2_1 U15994 ( .ip1(\pipeline/md/b [62]), .ip2(n21951), .op(n14749) );
  or2_1 U15995 ( .ip1(\pipeline/md/a [61]), .ip2(n14749), .op(n14751) );
  inv_1 U15996 ( .ip(\pipeline/md/b [61]), .op(n22744) );
  or2_1 U15997 ( .ip1(n22744), .ip2(n14749), .op(n14750) );
  nand2_1 U15998 ( .ip1(n14751), .ip2(n14750), .op(n14761) );
  inv_1 U15999 ( .ip(\pipeline/md/b [60]), .op(n22734) );
  nand2_1 U16000 ( .ip1(\pipeline/md/a [60]), .ip2(n22734), .op(n14755) );
  inv_1 U16001 ( .ip(\pipeline/md/b [58]), .op(n21308) );
  nand2_1 U16002 ( .ip1(\pipeline/md/a [58]), .ip2(n21308), .op(n21936) );
  inv_1 U16003 ( .ip(\pipeline/md/a [59]), .op(n14752) );
  nor2_1 U16004 ( .ip1(\pipeline/md/b [59]), .ip2(n14752), .op(n21935) );
  inv_1 U16005 ( .ip(n21935), .op(n21727) );
  nand4_1 U16006 ( .ip1(n14761), .ip2(n14755), .ip3(n21936), .ip4(n21727), 
        .op(n14753) );
  nor2_1 U16007 ( .ip1(n14754), .ip2(n14753), .op(n14768) );
  inv_1 U16008 ( .ip(\pipeline/md/a [60]), .op(n21735) );
  nor2_1 U16009 ( .ip1(\pipeline/md/a [61]), .ip2(n22744), .op(n14760) );
  inv_1 U16010 ( .ip(n14755), .op(n14758) );
  nor2_1 U16011 ( .ip1(\pipeline/md/a [58]), .ip2(n21308), .op(n21940) );
  inv_1 U16012 ( .ip(\pipeline/md/b [59]), .op(n14756) );
  nor2_1 U16013 ( .ip1(\pipeline/md/a [59]), .ip2(n14756), .op(n21934) );
  nor2_1 U16014 ( .ip1(n21940), .ip2(n21934), .op(n14757) );
  or2_1 U16015 ( .ip1(n21935), .ip2(n14757), .op(n21729) );
  nor2_1 U16016 ( .ip1(n14758), .ip2(n21729), .op(n14759) );
  not_ab_or_c_or_d U16017 ( .ip1(\pipeline/md/b [60]), .ip2(n21735), .ip3(
        n14760), .ip4(n14759), .op(n14763) );
  inv_1 U16018 ( .ip(n14761), .op(n14762) );
  nor2_1 U16019 ( .ip1(n14763), .ip2(n14762), .op(n14767) );
  inv_1 U16020 ( .ip(\pipeline/md/b [62]), .op(n21681) );
  nor2_1 U16021 ( .ip1(\pipeline/md/a [62]), .ip2(n21681), .op(n14766) );
  inv_1 U16022 ( .ip(\pipeline/md/state [0]), .op(n14764) );
  nor2_1 U16023 ( .ip1(\pipeline/md/state [1]), .ip2(n14764), .op(n14765) );
  inv_1 U16024 ( .ip(n14765), .op(n22665) );
  or2_1 U16025 ( .ip1(\pipeline/md/op [0]), .ip2(\pipeline/md/op [1]), .op(
        n15116) );
  nand2_1 U16026 ( .ip1(n14765), .ip2(n15116), .op(n14855) );
  or4_1 U16027 ( .ip1(n14768), .ip2(n14767), .ip3(n14766), .ip4(n14855), .op(
        n14769) );
  nand2_1 U16028 ( .ip1(n21683), .ip2(n14769), .op(n14770) );
  inv_1 U16029 ( .ip(n14770), .op(n21947) );
  nand2_1 U16030 ( .ip1(n14770), .ip2(n14771), .op(n21499) );
  inv_1 U16031 ( .ip(n21499), .op(n21649) );
  nand2_1 U16032 ( .ip1(n21649), .ip2(n20483), .op(n20649) );
  nand2_1 U16033 ( .ip1(n16237), .ip2(n14772), .op(n14773) );
  nand2_1 U16034 ( .ip1(n21649), .ip2(n14773), .op(n14774) );
  nand2_1 U16035 ( .ip1(n20649), .ip2(n14774), .op(n14775) );
  nand2_1 U16036 ( .ip1(n20645), .ip2(n14775), .op(n14816) );
  inv_1 U16037 ( .ip(n14776), .op(n14779) );
  nand2_1 U16038 ( .ip1(n14777), .ip2(n20431), .op(n14778) );
  nand2_1 U16039 ( .ip1(n14779), .ip2(n14778), .op(n18151) );
  nor2_1 U16040 ( .ip1(n14780), .ip2(n18151), .op(n14781) );
  nor2_1 U16041 ( .ip1(n14782), .ip2(n14781), .op(n20011) );
  nand2_1 U16042 ( .ip1(n20011), .ip2(n14783), .op(n14784) );
  nand2_1 U16043 ( .ip1(n14785), .ip2(n14784), .op(n20443) );
  nand2_1 U16044 ( .ip1(n14786), .ip2(n20443), .op(n20565) );
  nand2_1 U16045 ( .ip1(n14787), .ip2(n20565), .op(n14789) );
  nand2_1 U16046 ( .ip1(n14789), .ip2(n14788), .op(n20576) );
  nor2_1 U16047 ( .ip1(n14790), .ip2(n20576), .op(n14791) );
  nor2_1 U16048 ( .ip1(n14792), .ip2(n14791), .op(n20591) );
  nor2_1 U16049 ( .ip1(n20591), .ip2(n14793), .op(n20282) );
  nor2_1 U16050 ( .ip1(n20282), .ip2(n14794), .op(n14796) );
  nor2_1 U16051 ( .ip1(n14796), .ip2(n14795), .op(n20616) );
  inv_1 U16052 ( .ip(n20616), .op(n14798) );
  nand2_1 U16053 ( .ip1(n14798), .ip2(n14797), .op(n14799) );
  nand2_1 U16054 ( .ip1(n14800), .ip2(n14799), .op(n20151) );
  nor2_1 U16055 ( .ip1(\pipeline/md/b [25]), .ip2(n20151), .op(n14801) );
  or2_1 U16056 ( .ip1(\pipeline/md/a [25]), .ip2(n14801), .op(n20146) );
  nand2_1 U16057 ( .ip1(\pipeline/md/b [25]), .ip2(n20151), .op(n20149) );
  nand2_1 U16058 ( .ip1(n20146), .ip2(n20149), .op(n20626) );
  nand2_1 U16059 ( .ip1(n20626), .ip2(n14802), .op(n14803) );
  nand2_1 U16060 ( .ip1(n14804), .ip2(n14803), .op(n14806) );
  nor2_1 U16061 ( .ip1(\pipeline/md/b [27]), .ip2(n14806), .op(n14805) );
  nor2_1 U16062 ( .ip1(\pipeline/md/a [27]), .ip2(n14805), .op(n20639) );
  and2_1 U16063 ( .ip1(n14770), .ip2(n14765), .op(n21944) );
  inv_1 U16064 ( .ip(n14806), .op(n14809) );
  nor2_1 U16065 ( .ip1(n14809), .ip2(n15279), .op(n20638) );
  inv_1 U16066 ( .ip(n20638), .op(n14807) );
  nand3_1 U16067 ( .ip1(n20639), .ip2(n21944), .ip3(n14807), .op(n14815) );
  nand2_1 U16068 ( .ip1(n21947), .ip2(\pipeline/md/a [27]), .op(n14814) );
  inv_1 U16069 ( .ip(n22665), .op(n21440) );
  nand2_1 U16070 ( .ip1(n20638), .ip2(\pipeline/md/a [27]), .op(n14811) );
  nand2_1 U16071 ( .ip1(n14809), .ip2(n14808), .op(n14810) );
  nand2_1 U16072 ( .ip1(n14811), .ip2(n14810), .op(n14812) );
  nand2_1 U16073 ( .ip1(n21440), .ip2(n14812), .op(n14813) );
  nand4_1 U16074 ( .ip1(n14816), .ip2(n14815), .ip3(n14814), .ip4(n14813), 
        .op(n8419) );
  inv_1 U16075 ( .ip(\pipeline/md/state [1]), .op(n14817) );
  nor2_1 U16076 ( .ip1(\pipeline/md/state [0]), .ip2(n14817), .op(n20552) );
  inv_1 U16077 ( .ip(\pipeline/md_resp_result [31]), .op(n14819) );
  inv_1 U16078 ( .ip(\pipeline/md/a [31]), .op(n14818) );
  inv_1 U16079 ( .ip(\pipeline/md/out_sel [1]), .op(n14845) );
  nor2_1 U16080 ( .ip1(\pipeline/md/out_sel [0]), .ip2(n14845), .op(n14833) );
  mux2_1 U16081 ( .ip1(n14819), .ip2(n14818), .s(n14833), .op(n21666) );
  mux2_1 U16082 ( .ip1(\pipeline/md_resp_result [30]), .ip2(
        \pipeline/md/a [30]), .s(n14833), .op(n18855) );
  inv_1 U16083 ( .ip(\pipeline/md_resp_result [29]), .op(n14821) );
  mux2_1 U16084 ( .ip1(n14821), .ip2(n14820), .s(n14833), .op(n20664) );
  mux2_1 U16085 ( .ip1(\pipeline/md_resp_result [28]), .ip2(
        \pipeline/md/a [28]), .s(n14833), .op(n19016) );
  inv_1 U16086 ( .ip(\pipeline/md_resp_result [27]), .op(n14823) );
  buf_1 U16087 ( .ip(n14833), .op(n14842) );
  mux2_1 U16088 ( .ip1(n14823), .ip2(n14822), .s(n14842), .op(n15264) );
  mux2_1 U16089 ( .ip1(\pipeline/md_resp_result [26]), .ip2(
        \pipeline/md/a [26]), .s(n14833), .op(n20295) );
  mux2_1 U16090 ( .ip1(\pipeline/md_resp_result [22]), .ip2(
        \pipeline/md/a [22]), .s(n14833), .op(n18122) );
  mux2_1 U16091 ( .ip1(\pipeline/md_resp_result [23]), .ip2(
        \pipeline/md/a [23]), .s(n14842), .op(n18120) );
  mux2_1 U16092 ( .ip1(\pipeline/md_resp_result [21]), .ip2(
        \pipeline/md/a [21]), .s(n14842), .op(n20452) );
  mux2_1 U16093 ( .ip1(\pipeline/md_resp_result [19]), .ip2(
        \pipeline/md/a [19]), .s(n14833), .op(n20544) );
  inv_1 U16094 ( .ip(\pipeline/md_resp_result [18]), .op(n14825) );
  mux2_1 U16095 ( .ip1(n14825), .ip2(n14824), .s(n14842), .op(n20543) );
  inv_1 U16096 ( .ip(n20543), .op(n15205) );
  mux2_1 U16097 ( .ip1(\pipeline/md_resp_result [17]), .ip2(
        \pipeline/md/a [17]), .s(n14842), .op(n15178) );
  inv_1 U16098 ( .ip(\pipeline/md_resp_result [16]), .op(n18193) );
  mux2_1 U16099 ( .ip1(n18193), .ip2(n14826), .s(n14842), .op(n18184) );
  mux2_1 U16100 ( .ip1(\pipeline/md_resp_result [15]), .ip2(
        \pipeline/md/a [15]), .s(n14842), .op(n15153) );
  inv_1 U16101 ( .ip(\pipeline/md_resp_result [12]), .op(n15111) );
  mux2_1 U16102 ( .ip1(n15111), .ip2(n14868), .s(n14833), .op(n15102) );
  inv_1 U16103 ( .ip(n15102), .op(n14836) );
  inv_1 U16104 ( .ip(\pipeline/md_resp_result [11]), .op(n18065) );
  inv_1 U16105 ( .ip(\pipeline/md/a [11]), .op(n14827) );
  mux2_1 U16106 ( .ip1(n18065), .ip2(n14827), .s(n14842), .op(n18082) );
  inv_1 U16107 ( .ip(\pipeline/md_resp_result [10]), .op(n15083) );
  inv_1 U16108 ( .ip(\pipeline/md/a [10]), .op(n14828) );
  mux2_1 U16109 ( .ip1(n15083), .ip2(n14828), .s(n14833), .op(n18075) );
  mux2_1 U16110 ( .ip1(\pipeline/md_resp_result [9]), .ip2(\pipeline/md/a [9]), 
        .s(n14842), .op(n15049) );
  inv_1 U16111 ( .ip(\pipeline/md_resp_result [8]), .op(n18217) );
  mux2_1 U16112 ( .ip1(n18217), .ip2(n14829), .s(n14842), .op(n18208) );
  mux2_1 U16113 ( .ip1(\pipeline/md_resp_result [7]), .ip2(\pipeline/md/a [7]), 
        .s(n14842), .op(n15024) );
  inv_1 U16114 ( .ip(\pipeline/md_resp_result [6]), .op(n14830) );
  mux2_1 U16115 ( .ip1(n14830), .ip2(n14873), .s(n14833), .op(n14990) );
  mux2_1 U16116 ( .ip1(\pipeline/md_resp_result [5]), .ip2(\pipeline/md/a [5]), 
        .s(n14833), .op(n14976) );
  inv_1 U16117 ( .ip(\pipeline/md_resp_result [4]), .op(n14962) );
  inv_1 U16118 ( .ip(\pipeline/md/a [4]), .op(n14831) );
  mux2_1 U16119 ( .ip1(n14962), .ip2(n14831), .s(n14833), .op(n14945) );
  mux2_1 U16120 ( .ip1(\pipeline/md_resp_result [3]), .ip2(\pipeline/md/a [3]), 
        .s(n14842), .op(n17869) );
  mux2_1 U16121 ( .ip1(\pipeline/md_resp_result [1]), .ip2(\pipeline/md/a [1]), 
        .s(n14833), .op(n21256) );
  inv_1 U16122 ( .ip(n21256), .op(n14834) );
  inv_1 U16123 ( .ip(\pipeline/md_resp_result [0]), .op(n21523) );
  mux2_1 U16124 ( .ip1(n21523), .ip2(n14832), .s(n14833), .op(n21255) );
  inv_1 U16125 ( .ip(\pipeline/md/a [2]), .op(n17342) );
  mux2_1 U16126 ( .ip1(n14920), .ip2(n17342), .s(n14833), .op(n14849) );
  nand3_1 U16127 ( .ip1(n14834), .ip2(n21255), .ip3(n14849), .op(n17866) );
  nor2_1 U16128 ( .ip1(n17869), .ip2(n17866), .op(n14947) );
  nand2_1 U16129 ( .ip1(n14945), .ip2(n14947), .op(n14973) );
  nor2_1 U16130 ( .ip1(n14976), .ip2(n14973), .op(n14988) );
  nand2_1 U16131 ( .ip1(n14990), .ip2(n14988), .op(n15021) );
  nor2_1 U16132 ( .ip1(n15024), .ip2(n15021), .op(n18205) );
  nand2_1 U16133 ( .ip1(n18208), .ip2(n18205), .op(n15046) );
  nor2_1 U16134 ( .ip1(n15049), .ip2(n15046), .op(n18074) );
  nand2_1 U16135 ( .ip1(n18075), .ip2(n18074), .op(n18083) );
  inv_1 U16136 ( .ip(n18083), .op(n14835) );
  nand2_1 U16137 ( .ip1(n18082), .ip2(n14835), .op(n15099) );
  nor2_1 U16138 ( .ip1(n14836), .ip2(n15099), .op(n15121) );
  mux2_1 U16139 ( .ip1(\pipeline/md_resp_result [13]), .ip2(
        \pipeline/md/a [13]), .s(n14842), .op(n18157) );
  inv_1 U16140 ( .ip(n18157), .op(n14838) );
  inv_1 U16141 ( .ip(\pipeline/md_resp_result [14]), .op(n15142) );
  inv_1 U16142 ( .ip(\pipeline/md/a [14]), .op(n14837) );
  mux2_1 U16143 ( .ip1(n15142), .ip2(n14837), .s(n14842), .op(n18162) );
  nand3_1 U16144 ( .ip1(n15121), .ip2(n14838), .ip3(n18162), .op(n15150) );
  nor2_1 U16145 ( .ip1(n15153), .ip2(n15150), .op(n18182) );
  nand2_1 U16146 ( .ip1(n18184), .ip2(n18182), .op(n15175) );
  nor2_1 U16147 ( .ip1(n15178), .ip2(n15175), .op(n15199) );
  inv_1 U16148 ( .ip(n15199), .op(n14839) );
  nor2_1 U16149 ( .ip1(n15205), .ip2(n14839), .op(n20537) );
  inv_1 U16150 ( .ip(n20537), .op(n14840) );
  nor2_1 U16151 ( .ip1(n20544), .ip2(n14840), .op(n18251) );
  inv_1 U16152 ( .ip(\pipeline/md_resp_result [20]), .op(n14841) );
  mux2_1 U16153 ( .ip1(n14841), .ip2(n14885), .s(n14842), .op(n18253) );
  nand2_1 U16154 ( .ip1(n18251), .ip2(n18253), .op(n20449) );
  nor2_1 U16155 ( .ip1(n20452), .ip2(n20449), .op(n18101) );
  inv_1 U16156 ( .ip(n18101), .op(n18121) );
  nor3_1 U16157 ( .ip1(n18122), .ip2(n18120), .ip3(n18121), .op(n21958) );
  mux2_1 U16158 ( .ip1(\pipeline/md_resp_result [24]), .ip2(
        \pipeline/md/a [24]), .s(n14842), .op(n21959) );
  inv_1 U16159 ( .ip(n21959), .op(n14844) );
  inv_1 U16160 ( .ip(\pipeline/md_resp_result [25]), .op(n14843) );
  inv_1 U16161 ( .ip(\pipeline/md/a [25]), .op(n20148) );
  mux2_1 U16162 ( .ip1(n14843), .ip2(n20148), .s(n14842), .op(n15220) );
  nand3_1 U16163 ( .ip1(n21958), .ip2(n14844), .ip3(n15220), .op(n20292) );
  nor2_1 U16164 ( .ip1(n20295), .ip2(n20292), .op(n15262) );
  nand2_1 U16165 ( .ip1(n15264), .ip2(n15262), .op(n19013) );
  nor2_1 U16166 ( .ip1(n19016), .ip2(n19013), .op(n20666) );
  nand2_1 U16167 ( .ip1(n20664), .ip2(n20666), .op(n18852) );
  nor2_1 U16168 ( .ip1(n18855), .ip2(n18852), .op(n21658) );
  and2_1 U16169 ( .ip1(n21666), .ip2(n21658), .op(n21506) );
  inv_1 U16170 ( .ip(\pipeline/md/result [32]), .op(n21510) );
  nand2_1 U16171 ( .ip1(n21506), .ip2(n21510), .op(n21263) );
  or2_1 U16172 ( .ip1(\pipeline/md/result [33]), .ip2(n21263), .op(n14846) );
  nor2_1 U16173 ( .ip1(n14846), .ip2(\pipeline/md/result [34]), .op(n17873) );
  nand2_1 U16174 ( .ip1(\pipeline/md/out_sel [0]), .ip2(n14845), .op(n21662)
         );
  inv_1 U16175 ( .ip(n21662), .op(n21960) );
  nand2_1 U16176 ( .ip1(\pipeline/md/negate_output ), .ip2(n21960), .op(n21505) );
  not_ab_or_c_or_d U16177 ( .ip1(\pipeline/md/result [34]), .ip2(n14846), 
        .ip3(n17873), .ip4(n21505), .op(n14853) );
  inv_1 U16178 ( .ip(n21255), .op(n21520) );
  nor2_1 U16179 ( .ip1(n21256), .ip2(n21520), .op(n14847) );
  inv_1 U16180 ( .ip(\pipeline/md/negate_output ), .op(n21659) );
  nor2_1 U16181 ( .ip1(n14847), .ip2(n21659), .op(n14848) );
  xor2_1 U16182 ( .ip1(n14849), .ip2(n14848), .op(n14850) );
  inv_1 U16183 ( .ip(n20552), .op(n21967) );
  nor2_1 U16184 ( .ip1(n21960), .ip2(n21967), .op(n21972) );
  inv_1 U16185 ( .ip(n21972), .op(n15265) );
  nor2_1 U16186 ( .ip1(n14850), .ip2(n15265), .op(n14852) );
  or2_1 U16187 ( .ip1(\pipeline/md/negate_output ), .ip2(n21662), .op(n15200)
         );
  inv_1 U16188 ( .ip(n15200), .op(n21509) );
  nand2_1 U16189 ( .ip1(n20552), .ip2(n21509), .op(n15267) );
  inv_1 U16190 ( .ip(\pipeline/md/result [34]), .op(n22510) );
  nor2_1 U16191 ( .ip1(n15267), .ip2(n22510), .op(n14851) );
  not_ab_or_c_or_d U16192 ( .ip1(n20552), .ip2(n14853), .ip3(n14852), .ip4(
        n14851), .op(n14928) );
  inv_1 U16193 ( .ip(\pipeline/md/counter [1]), .op(n14854) );
  nor2_1 U16194 ( .ip1(\pipeline/md/counter [0]), .ip2(n14854), .op(n15188) );
  inv_1 U16195 ( .ip(n14855), .op(n18216) );
  inv_1 U16196 ( .ip(\pipeline/md/counter [4]), .op(n14911) );
  nand2_1 U16197 ( .ip1(n18216), .ip2(n14911), .op(n21515) );
  nor2_1 U16198 ( .ip1(\pipeline/md/counter [2]), .ip2(
        \pipeline/md/counter [3]), .op(n14914) );
  inv_1 U16199 ( .ip(\pipeline/md/counter [0]), .op(n14856) );
  or2_1 U16200 ( .ip1(\pipeline/md/counter [1]), .ip2(n14856), .op(n14972) );
  nor2_1 U16201 ( .ip1(n14857), .ip2(n14972), .op(n14858) );
  inv_1 U16202 ( .ip(\pipeline/md/counter [3]), .op(n14943) );
  not_ab_or_c_or_d U16203 ( .ip1(\pipeline/md/a [10]), .ip2(n15188), .ip3(
        n14858), .ip4(n14943), .op(n14861) );
  nand2_1 U16204 ( .ip1(\pipeline/md/counter [0]), .ip2(
        \pipeline/md/counter [1]), .op(n15289) );
  inv_1 U16205 ( .ip(n15289), .op(n20554) );
  nand2_1 U16206 ( .ip1(\pipeline/md/a [11]), .ip2(n20554), .op(n14860) );
  nor2_1 U16207 ( .ip1(\pipeline/md/counter [0]), .ip2(
        \pipeline/md/counter [1]), .op(n17747) );
  nand2_1 U16208 ( .ip1(\pipeline/md/a [8]), .ip2(n17747), .op(n14859) );
  nand3_1 U16209 ( .ip1(n14861), .ip2(n14860), .ip3(n14859), .op(n14867) );
  inv_1 U16210 ( .ip(n14972), .op(n21272) );
  inv_1 U16211 ( .ip(n15188), .op(n15006) );
  nor2_1 U16212 ( .ip1(n15006), .ip2(n17342), .op(n14862) );
  not_ab_or_c_or_d U16213 ( .ip1(n21272), .ip2(\pipeline/md/a [1]), .ip3(
        \pipeline/md/counter [3]), .ip4(n14862), .op(n14865) );
  nand2_1 U16214 ( .ip1(n20554), .ip2(\pipeline/md/a [3]), .op(n14864) );
  nand2_1 U16215 ( .ip1(n17747), .ip2(\pipeline/md/a [0]), .op(n14863) );
  nand3_1 U16216 ( .ip1(n14865), .ip2(n14864), .ip3(n14863), .op(n14866) );
  nand2_1 U16217 ( .ip1(n14867), .ip2(n14866), .op(n14881) );
  inv_1 U16218 ( .ip(n17747), .op(n18213) );
  nor2_1 U16219 ( .ip1(n14868), .ip2(n18213), .op(n14872) );
  nand2_1 U16220 ( .ip1(\pipeline/md/a [13]), .ip2(n21272), .op(n14870) );
  nand2_1 U16221 ( .ip1(\pipeline/md/a [14]), .ip2(n15188), .op(n14869) );
  nand3_1 U16222 ( .ip1(\pipeline/md/counter [3]), .ip2(n14870), .ip3(n14869), 
        .op(n14871) );
  not_ab_or_c_or_d U16223 ( .ip1(n20554), .ip2(\pipeline/md/a [15]), .ip3(
        n14872), .ip4(n14871), .op(n14879) );
  nor2_1 U16224 ( .ip1(n14873), .ip2(n15006), .op(n14877) );
  nand2_1 U16225 ( .ip1(\pipeline/md/a [7]), .ip2(n20554), .op(n14875) );
  nand2_1 U16226 ( .ip1(\pipeline/md/a [4]), .ip2(n17747), .op(n14874) );
  nand3_1 U16227 ( .ip1(n14943), .ip2(n14875), .ip3(n14874), .op(n14876) );
  not_ab_or_c_or_d U16228 ( .ip1(n21272), .ip2(\pipeline/md/a [5]), .ip3(
        n14877), .ip4(n14876), .op(n14878) );
  or2_1 U16229 ( .ip1(n14879), .ip2(n14878), .op(n14880) );
  mux2_1 U16230 ( .ip1(n14881), .ip2(n14880), .s(\pipeline/md/counter [2]), 
        .op(n14910) );
  nand2_1 U16231 ( .ip1(n20554), .ip2(\pipeline/md/a [19]), .op(n14884) );
  nand2_1 U16232 ( .ip1(\pipeline/md/a [17]), .ip2(n21272), .op(n14883) );
  nand2_1 U16233 ( .ip1(\pipeline/md/a [18]), .ip2(n15188), .op(n14882) );
  nand3_1 U16234 ( .ip1(n14884), .ip2(n14883), .ip3(n14882), .op(n14908) );
  nor2_1 U16235 ( .ip1(n14885), .ip2(n18213), .op(n14889) );
  nor2_1 U16236 ( .ip1(n14886), .ip2(n15006), .op(n14887) );
  ab_or_c_or_d U16237 ( .ip1(n21272), .ip2(\pipeline/md/a [21]), .ip3(
        \pipeline/md/counter [3]), .ip4(n14887), .op(n14888) );
  not_ab_or_c_or_d U16238 ( .ip1(n20554), .ip2(\pipeline/md/a [23]), .ip3(
        n14889), .ip4(n14888), .op(n14897) );
  nor2_1 U16239 ( .ip1(n14890), .ip2(n15006), .op(n14894) );
  nand2_1 U16240 ( .ip1(\pipeline/md/a [29]), .ip2(n21272), .op(n14892) );
  nand2_1 U16241 ( .ip1(\pipeline/md/a [28]), .ip2(n17747), .op(n14891) );
  nand3_1 U16242 ( .ip1(\pipeline/md/counter [3]), .ip2(n14892), .ip3(n14891), 
        .op(n14893) );
  not_ab_or_c_or_d U16243 ( .ip1(n20554), .ip2(\pipeline/md/a [31]), .ip3(
        n14894), .ip4(n14893), .op(n14896) );
  inv_1 U16244 ( .ip(\pipeline/md/counter [2]), .op(n14895) );
  nor3_1 U16245 ( .ip1(n14897), .ip2(n14896), .ip3(n14895), .op(n14907) );
  nor2_1 U16246 ( .ip1(\pipeline/md/counter [2]), .ip2(n14943), .op(n17760) );
  nand2_1 U16247 ( .ip1(\pipeline/md/a [27]), .ip2(n20554), .op(n14901) );
  nand2_1 U16248 ( .ip1(\pipeline/md/a [24]), .ip2(n17747), .op(n14900) );
  nand2_1 U16249 ( .ip1(\pipeline/md/a [25]), .ip2(n21272), .op(n14899) );
  nand2_1 U16250 ( .ip1(\pipeline/md/a [26]), .ip2(n15188), .op(n14898) );
  nand4_1 U16251 ( .ip1(n14901), .ip2(n14900), .ip3(n14899), .ip4(n14898), 
        .op(n14902) );
  nand2_1 U16252 ( .ip1(n17760), .ip2(n14902), .op(n14905) );
  inv_1 U16253 ( .ip(n14914), .op(n14903) );
  nor2_1 U16254 ( .ip1(n18213), .ip2(n14903), .op(n17751) );
  nand2_1 U16255 ( .ip1(\pipeline/md/a [16]), .ip2(n17751), .op(n14904) );
  nand3_1 U16256 ( .ip1(\pipeline/md/counter [4]), .ip2(n14905), .ip3(n14904), 
        .op(n14906) );
  not_ab_or_c_or_d U16257 ( .ip1(n14914), .ip2(n14908), .ip3(n14907), .ip4(
        n14906), .op(n14909) );
  inv_1 U16258 ( .ip(n15116), .op(n21248) );
  nand2_1 U16259 ( .ip1(n21248), .ip2(n21440), .op(n18219) );
  not_ab_or_c_or_d U16260 ( .ip1(n14911), .ip2(n14910), .ip3(n14909), .ip4(
        n18219), .op(n14912) );
  or2_1 U16261 ( .ip1(n14912), .ip2(n20552), .op(n14913) );
  nor2_1 U16262 ( .ip1(n14913), .ip2(n14770), .op(n21517) );
  inv_1 U16263 ( .ip(n21517), .op(n21250) );
  nand2_1 U16264 ( .ip1(n14914), .ip2(n21250), .op(n15163) );
  nor2_1 U16265 ( .ip1(n21515), .ip2(n15163), .op(n21271) );
  nand2_1 U16266 ( .ip1(n15188), .ip2(n21271), .op(n14927) );
  nor2_1 U16267 ( .ip1(n22665), .ip2(n21517), .op(n21251) );
  inv_1 U16268 ( .ip(\pipeline/md_resp_result [1]), .op(n14916) );
  and2_1 U16269 ( .ip1(\pipeline/md_resp_result [0]), .ip2(\pipeline/md/b [0]), 
        .op(n14915) );
  nor2_1 U16270 ( .ip1(\pipeline/md/b [1]), .ip2(n14915), .op(n21245) );
  or2_1 U16271 ( .ip1(n14916), .ip2(n21245), .op(n14917) );
  nand3_1 U16272 ( .ip1(\pipeline/md/b [1]), .ip2(\pipeline/md_resp_result [0]), .ip3(\pipeline/md/b [0]), .op(n21247) );
  nand2_1 U16273 ( .ip1(n14917), .ip2(n21247), .op(n14918) );
  nor2_1 U16274 ( .ip1(n14918), .ip2(\pipeline/md/b [2]), .op(n14931) );
  inv_1 U16275 ( .ip(n14918), .op(n14919) );
  nor2_1 U16276 ( .ip1(n14919), .ip2(n17341), .op(n14929) );
  nor3_1 U16277 ( .ip1(n14931), .ip2(n14929), .ip3(n15116), .op(n14921) );
  nand3_1 U16278 ( .ip1(n21251), .ip2(n14921), .ip3(n14920), .op(n14926) );
  inv_1 U16279 ( .ip(n14921), .op(n14922) );
  nand2_1 U16280 ( .ip1(n14765), .ip2(n14922), .op(n14923) );
  nand2_1 U16281 ( .ip1(n21250), .ip2(n14923), .op(n14924) );
  nand2_1 U16282 ( .ip1(\pipeline/md_resp_result [2]), .ip2(n14924), .op(
        n14925) );
  nand4_1 U16283 ( .ip1(n14928), .ip2(n14927), .ip3(n14926), .ip4(n14925), 
        .op(n8632) );
  nor2_1 U16284 ( .ip1(\pipeline/md_resp_result [2]), .ip2(n14929), .op(n14932) );
  nor2_1 U16285 ( .ip1(n14931), .ip2(n14932), .op(n14930) );
  nor2_1 U16286 ( .ip1(\pipeline/md/b [3]), .ip2(n14930), .op(n17865) );
  inv_1 U16287 ( .ip(n17865), .op(n17861) );
  inv_1 U16288 ( .ip(\pipeline/md_resp_result [3]), .op(n14935) );
  inv_1 U16289 ( .ip(n14931), .op(n14934) );
  inv_1 U16290 ( .ip(n14932), .op(n14933) );
  nand3_1 U16291 ( .ip1(\pipeline/md/b [3]), .ip2(n14934), .ip3(n14933), .op(
        n17860) );
  nand2_1 U16292 ( .ip1(n14935), .ip2(n17860), .op(n17864) );
  nand2_1 U16293 ( .ip1(n17861), .ip2(n17864), .op(n14937) );
  nand2_1 U16294 ( .ip1(n14936), .ip2(n14937), .op(n14964) );
  inv_1 U16295 ( .ip(n14937), .op(n14938) );
  nand2_1 U16296 ( .ip1(\pipeline/md/b [4]), .ip2(n14938), .op(n14961) );
  nand3_1 U16297 ( .ip1(n21248), .ip2(n14964), .ip3(n14961), .op(n14940) );
  nor2_1 U16298 ( .ip1(\pipeline/md_resp_result [4]), .ip2(n14940), .op(n14939) );
  nand2_1 U16299 ( .ip1(n21251), .ip2(n14939), .op(n14960) );
  nand2_1 U16300 ( .ip1(n14765), .ip2(n14940), .op(n14941) );
  nand2_1 U16301 ( .ip1(n21250), .ip2(n14941), .op(n14942) );
  nand2_1 U16302 ( .ip1(n14942), .ip2(\pipeline/md_resp_result [4]), .op(
        n14959) );
  nor2_1 U16303 ( .ip1(n18213), .ip2(n21517), .op(n21977) );
  nand2_1 U16304 ( .ip1(\pipeline/md/counter [2]), .ip2(n14943), .op(n18098)
         );
  nor2_1 U16305 ( .ip1(n21515), .ip2(n18098), .op(n15020) );
  nand2_1 U16306 ( .ip1(n21977), .ip2(n15020), .op(n14958) );
  nor2_1 U16307 ( .ip1(n14947), .ip2(n21659), .op(n14944) );
  nor2_1 U16308 ( .ip1(n14945), .ip2(n14944), .op(n14951) );
  or2_1 U16309 ( .ip1(\pipeline/md/negate_output ), .ip2(n21960), .op(n18073)
         );
  inv_1 U16310 ( .ip(n18073), .op(n20669) );
  inv_1 U16311 ( .ip(n14945), .op(n14946) );
  nor2_1 U16312 ( .ip1(n14947), .ip2(n14946), .op(n14948) );
  nor2_1 U16313 ( .ip1(n21960), .ip2(n14948), .op(n14949) );
  nor2_1 U16314 ( .ip1(n20669), .ip2(n14949), .op(n14950) );
  nor2_1 U16315 ( .ip1(n14951), .ip2(n14950), .op(n14956) );
  inv_1 U16316 ( .ip(n17873), .op(n17872) );
  nor2_1 U16317 ( .ip1(\pipeline/md/result [35]), .ip2(n17872), .op(n14977) );
  nor2_1 U16318 ( .ip1(n21967), .ip2(n21659), .op(n17871) );
  inv_1 U16319 ( .ip(n17871), .op(n21966) );
  nor3_1 U16320 ( .ip1(\pipeline/md/result [36]), .ip2(n14977), .ip3(n21966), 
        .op(n14954) );
  inv_1 U16321 ( .ip(n14977), .op(n14952) );
  inv_1 U16322 ( .ip(\pipeline/md/result [36]), .op(n22526) );
  not_ab_or_c_or_d U16323 ( .ip1(\pipeline/md/negate_output ), .ip2(n14952), 
        .ip3(n22526), .ip4(n21967), .op(n14953) );
  nor3_1 U16324 ( .ip1(n21972), .ip2(n14954), .ip3(n14953), .op(n14955) );
  or2_1 U16325 ( .ip1(n14956), .ip2(n14955), .op(n14957) );
  nand4_1 U16326 ( .ip1(n14960), .ip2(n14959), .ip3(n14958), .ip4(n14957), 
        .op(n8630) );
  nand2_1 U16327 ( .ip1(n14962), .ip2(n14961), .op(n14963) );
  nand2_1 U16328 ( .ip1(n14964), .ip2(n14963), .op(n14966) );
  nand2_1 U16329 ( .ip1(n14965), .ip2(n14966), .op(n15000) );
  inv_1 U16330 ( .ip(n14966), .op(n14967) );
  nand2_1 U16331 ( .ip1(\pipeline/md/b [5]), .ip2(n14967), .op(n14995) );
  nand3_1 U16332 ( .ip1(n21248), .ip2(n15000), .ip3(n14995), .op(n14969) );
  nor2_1 U16333 ( .ip1(\pipeline/md_resp_result [5]), .ip2(n14969), .op(n14968) );
  nand2_1 U16334 ( .ip1(n21251), .ip2(n14968), .op(n14985) );
  nand2_1 U16335 ( .ip1(n14765), .ip2(n14969), .op(n14970) );
  nand2_1 U16336 ( .ip1(n21250), .ip2(n14970), .op(n14971) );
  nand2_1 U16337 ( .ip1(n14971), .ip2(\pipeline/md_resp_result [5]), .op(
        n14984) );
  nor2_1 U16338 ( .ip1(n14972), .ip2(n21517), .op(n20680) );
  nand2_1 U16339 ( .ip1(n20680), .ip2(n15020), .op(n14983) );
  nand2_1 U16340 ( .ip1(\pipeline/md/negate_output ), .ip2(n14973), .op(n14975) );
  nor2_1 U16341 ( .ip1(n14976), .ip2(n14975), .op(n14974) );
  not_ab_or_c_or_d U16342 ( .ip1(n14976), .ip2(n14975), .ip3(n21960), .ip4(
        n14974), .op(n14981) );
  nand2_1 U16343 ( .ip1(n14977), .ip2(n22526), .op(n14986) );
  inv_1 U16344 ( .ip(\pipeline/md/result [37]), .op(n22542) );
  and3_1 U16345 ( .ip1(n17871), .ip2(n14986), .ip3(n22542), .op(n14979) );
  not_ab_or_c_or_d U16346 ( .ip1(\pipeline/md/negate_output ), .ip2(n14986), 
        .ip3(n22542), .ip4(n21967), .op(n14978) );
  nor3_1 U16347 ( .ip1(n21972), .ip2(n14979), .ip3(n14978), .op(n14980) );
  or2_1 U16348 ( .ip1(n14981), .ip2(n14980), .op(n14982) );
  nand4_1 U16349 ( .ip1(n14985), .ip2(n14984), .ip3(n14983), .ip4(n14982), 
        .op(n8629) );
  or2_1 U16350 ( .ip1(\pipeline/md/result [37]), .ip2(n14986), .op(n14987) );
  nor2_1 U16351 ( .ip1(n14987), .ip2(\pipeline/md/result [38]), .op(n15026) );
  not_ab_or_c_or_d U16352 ( .ip1(\pipeline/md/result [38]), .ip2(n14987), 
        .ip3(n15026), .ip4(n21505), .op(n14994) );
  nor2_1 U16353 ( .ip1(n14988), .ip2(n21659), .op(n14989) );
  xor2_1 U16354 ( .ip1(n14990), .ip2(n14989), .op(n14991) );
  nor2_1 U16355 ( .ip1(n14991), .ip2(n15265), .op(n14993) );
  inv_1 U16356 ( .ip(\pipeline/md/result [38]), .op(n22552) );
  nor2_1 U16357 ( .ip1(n22552), .ip2(n15267), .op(n14992) );
  not_ab_or_c_or_d U16358 ( .ip1(n20552), .ip2(n14994), .ip3(n14993), .ip4(
        n14992), .op(n15010) );
  nor2_1 U16359 ( .ip1(n18216), .ip2(n21517), .op(n22738) );
  inv_1 U16360 ( .ip(\pipeline/md/b [6]), .op(n14998) );
  inv_1 U16361 ( .ip(\pipeline/md_resp_result [5]), .op(n14996) );
  nand2_1 U16362 ( .ip1(n14996), .ip2(n14995), .op(n14999) );
  nand2_1 U16363 ( .ip1(n15000), .ip2(n14999), .op(n14997) );
  nand2_1 U16364 ( .ip1(n14998), .ip2(n14997), .op(n15011) );
  nand3_1 U16365 ( .ip1(\pipeline/md/b [6]), .ip2(n15000), .ip3(n14999), .op(
        n15004) );
  nand2_1 U16366 ( .ip1(n15011), .ip2(n15004), .op(n15001) );
  nand2_1 U16367 ( .ip1(n14765), .ip2(n15001), .op(n15002) );
  nand2_1 U16368 ( .ip1(n22738), .ip2(n15002), .op(n15003) );
  nand2_1 U16369 ( .ip1(\pipeline/md_resp_result [6]), .ip2(n15003), .op(
        n15009) );
  nor2_1 U16370 ( .ip1(n18219), .ip2(n21517), .op(n22750) );
  inv_1 U16371 ( .ip(n15004), .op(n15005) );
  nor2_1 U16372 ( .ip1(\pipeline/md_resp_result [6]), .ip2(n15005), .op(n15012) );
  nand3_1 U16373 ( .ip1(n22750), .ip2(n15012), .ip3(n15011), .op(n15008) );
  nor2_1 U16374 ( .ip1(n15006), .ip2(n21517), .op(n20306) );
  nand2_1 U16375 ( .ip1(n15020), .ip2(n20306), .op(n15007) );
  nand4_1 U16376 ( .ip1(n15010), .ip2(n15009), .ip3(n15008), .ip4(n15007), 
        .op(n8628) );
  inv_1 U16377 ( .ip(n15011), .op(n15013) );
  nor2_1 U16378 ( .ip1(n15013), .ip2(n15012), .op(n15014) );
  nand2_1 U16379 ( .ip1(\pipeline/md/b [7]), .ip2(n15014), .op(n15036) );
  nor2_1 U16380 ( .ip1(\pipeline/md/b [7]), .ip2(n15014), .op(n15034) );
  inv_1 U16381 ( .ip(n15034), .op(n15015) );
  nand3_1 U16382 ( .ip1(n21248), .ip2(n15036), .ip3(n15015), .op(n15017) );
  nor2_1 U16383 ( .ip1(\pipeline/md_resp_result [7]), .ip2(n15017), .op(n15016) );
  nand2_1 U16384 ( .ip1(n21251), .ip2(n15016), .op(n15033) );
  nand2_1 U16385 ( .ip1(n21440), .ip2(n15017), .op(n15018) );
  nand2_1 U16386 ( .ip1(n21250), .ip2(n15018), .op(n15019) );
  nand2_1 U16387 ( .ip1(n15019), .ip2(\pipeline/md_resp_result [7]), .op(
        n15032) );
  nor2_1 U16388 ( .ip1(n15289), .ip2(n21517), .op(n21671) );
  nand2_1 U16389 ( .ip1(n21671), .ip2(n15020), .op(n15031) );
  nand2_1 U16390 ( .ip1(\pipeline/md/negate_output ), .ip2(n15021), .op(n15023) );
  nor2_1 U16391 ( .ip1(n15024), .ip2(n15023), .op(n15022) );
  not_ab_or_c_or_d U16392 ( .ip1(n15024), .ip2(n15023), .ip3(n21960), .ip4(
        n15022), .op(n15029) );
  inv_1 U16393 ( .ip(n15026), .op(n15050) );
  inv_1 U16394 ( .ip(\pipeline/md/result [39]), .op(n22558) );
  nor2_1 U16395 ( .ip1(n21967), .ip2(n22558), .op(n15025) );
  not_ab_or_c_or_d U16396 ( .ip1(n17871), .ip2(n15050), .ip3(n21972), .ip4(
        n15025), .op(n15028) );
  nor3_1 U16397 ( .ip1(n22558), .ip2(n15026), .ip3(n21505), .op(n15027) );
  or3_1 U16398 ( .ip1(n15029), .ip2(n15028), .ip3(n15027), .op(n15030) );
  nand4_1 U16399 ( .ip1(n15033), .ip2(n15032), .ip3(n15031), .ip4(n15030), 
        .op(n8627) );
  inv_1 U16400 ( .ip(\pipeline/md_resp_result [7]), .op(n15035) );
  or2_1 U16401 ( .ip1(n15035), .ip2(n15034), .op(n15037) );
  nand2_1 U16402 ( .ip1(n15037), .ip2(n15036), .op(n15038) );
  nor2_1 U16403 ( .ip1(\pipeline/md/b [8]), .ip2(n15038), .op(n18221) );
  and2_1 U16404 ( .ip1(\pipeline/md/b [8]), .ip2(n15038), .op(n18220) );
  nor2_1 U16405 ( .ip1(\pipeline/md_resp_result [8]), .ip2(n18220), .op(n15039) );
  nor2_1 U16406 ( .ip1(n18221), .ip2(n15039), .op(n15040) );
  nand2_1 U16407 ( .ip1(\pipeline/md/b [9]), .ip2(n15040), .op(n15063) );
  inv_1 U16408 ( .ip(n15063), .op(n15041) );
  nor2_1 U16409 ( .ip1(\pipeline/md/b [9]), .ip2(n15040), .op(n15061) );
  or3_1 U16410 ( .ip1(n15041), .ip2(n15061), .ip3(n15116), .op(n15043) );
  nor2_1 U16411 ( .ip1(\pipeline/md_resp_result [9]), .ip2(n15043), .op(n15042) );
  nand2_1 U16412 ( .ip1(n21251), .ip2(n15042), .op(n15060) );
  inv_1 U16413 ( .ip(n22665), .op(n20310) );
  nand2_1 U16414 ( .ip1(n20310), .ip2(n15043), .op(n15044) );
  nand2_1 U16415 ( .ip1(n21250), .ip2(n15044), .op(n15045) );
  nand2_1 U16416 ( .ip1(n15045), .ip2(\pipeline/md_resp_result [9]), .op(
        n15059) );
  inv_1 U16417 ( .ip(n17760), .op(n15255) );
  nor2_1 U16418 ( .ip1(n15255), .ip2(n21515), .op(n18211) );
  nand2_1 U16419 ( .ip1(n20680), .ip2(n18211), .op(n15058) );
  nand2_1 U16420 ( .ip1(\pipeline/md/negate_output ), .ip2(n15046), .op(n15048) );
  nor2_1 U16421 ( .ip1(n15049), .ip2(n15048), .op(n15047) );
  not_ab_or_c_or_d U16422 ( .ip1(n15049), .ip2(n15048), .ip3(n21960), .ip4(
        n15047), .op(n15056) );
  nor2_1 U16423 ( .ip1(\pipeline/md/result [39]), .ip2(n15050), .op(n18202) );
  inv_1 U16424 ( .ip(\pipeline/md/result [40]), .op(n18204) );
  nand2_1 U16425 ( .ip1(n18202), .ip2(n18204), .op(n15071) );
  inv_1 U16426 ( .ip(n15071), .op(n15051) );
  nor3_1 U16427 ( .ip1(\pipeline/md/result [41]), .ip2(n21966), .ip3(n15051), 
        .op(n15054) );
  inv_1 U16428 ( .ip(\pipeline/md/result [41]), .op(n15052) );
  not_ab_or_c_or_d U16429 ( .ip1(\pipeline/md/negate_output ), .ip2(n15071), 
        .ip3(n15052), .ip4(n21967), .op(n15053) );
  nor3_1 U16430 ( .ip1(n21972), .ip2(n15054), .ip3(n15053), .op(n15055) );
  or2_1 U16431 ( .ip1(n15056), .ip2(n15055), .op(n15057) );
  nand4_1 U16432 ( .ip1(n15060), .ip2(n15059), .ip3(n15058), .ip4(n15057), 
        .op(n8625) );
  inv_1 U16433 ( .ip(\pipeline/md_resp_result [9]), .op(n15062) );
  or2_1 U16434 ( .ip1(n15062), .ip2(n15061), .op(n15064) );
  nand2_1 U16435 ( .ip1(n15064), .ip2(n15063), .op(n15065) );
  nand2_1 U16436 ( .ip1(\pipeline/md/b [10]), .ip2(n15065), .op(n15084) );
  nor2_1 U16437 ( .ip1(\pipeline/md/b [10]), .ip2(n15065), .op(n15082) );
  inv_1 U16438 ( .ip(n15082), .op(n15066) );
  nand3_1 U16439 ( .ip1(n21248), .ip2(n15084), .ip3(n15066), .op(n15068) );
  nor2_1 U16440 ( .ip1(\pipeline/md_resp_result [10]), .ip2(n15068), .op(
        n15067) );
  nand2_1 U16441 ( .ip1(n21251), .ip2(n15067), .op(n15081) );
  nand2_1 U16442 ( .ip1(n20310), .ip2(n15068), .op(n15069) );
  nand2_1 U16443 ( .ip1(n21250), .ip2(n15069), .op(n15070) );
  nand2_1 U16444 ( .ip1(n15070), .ip2(\pipeline/md_resp_result [10]), .op(
        n15080) );
  nand2_1 U16445 ( .ip1(n20306), .ip2(n18211), .op(n15079) );
  or2_1 U16446 ( .ip1(\pipeline/md/result [41]), .ip2(n15071), .op(n15072) );
  nor2_1 U16447 ( .ip1(n15072), .ip2(\pipeline/md/result [42]), .op(n15096) );
  not_ab_or_c_or_d U16448 ( .ip1(\pipeline/md/result [42]), .ip2(n15072), 
        .ip3(n15096), .ip4(n21505), .op(n15076) );
  or2_1 U16449 ( .ip1(n18074), .ip2(n21659), .op(n15074) );
  nor2_1 U16450 ( .ip1(n18075), .ip2(n15074), .op(n15073) );
  not_ab_or_c_or_d U16451 ( .ip1(n18075), .ip2(n15074), .ip3(n21960), .ip4(
        n15073), .op(n15075) );
  not_ab_or_c_or_d U16452 ( .ip1(\pipeline/md/result [42]), .ip2(n21509), 
        .ip3(n15076), .ip4(n15075), .op(n15077) );
  or2_1 U16453 ( .ip1(n15077), .ip2(n21967), .op(n15078) );
  nand4_1 U16454 ( .ip1(n15081), .ip2(n15080), .ip3(n15079), .ip4(n15078), 
        .op(n8624) );
  or2_1 U16455 ( .ip1(n15083), .ip2(n15082), .op(n15085) );
  nand2_1 U16456 ( .ip1(n15085), .ip2(n15084), .op(n15086) );
  nor2_1 U16457 ( .ip1(\pipeline/md/b [11]), .ip2(n15086), .op(n18068) );
  inv_1 U16458 ( .ip(n15086), .op(n15087) );
  nor2_1 U16459 ( .ip1(n15088), .ip2(n15087), .op(n18067) );
  nor2_1 U16460 ( .ip1(\pipeline/md_resp_result [11]), .ip2(n18067), .op(
        n15089) );
  nor2_1 U16461 ( .ip1(n18068), .ip2(n15089), .op(n15090) );
  nand2_1 U16462 ( .ip1(\pipeline/md/b [12]), .ip2(n15090), .op(n15112) );
  nor2_1 U16463 ( .ip1(\pipeline/md/b [12]), .ip2(n15090), .op(n15110) );
  inv_1 U16464 ( .ip(n15110), .op(n15091) );
  nand3_1 U16465 ( .ip1(n21248), .ip2(n15112), .ip3(n15091), .op(n15093) );
  nor2_1 U16466 ( .ip1(\pipeline/md_resp_result [12]), .ip2(n15093), .op(
        n15092) );
  nand2_1 U16467 ( .ip1(n21251), .ip2(n15092), .op(n15109) );
  nand2_1 U16468 ( .ip1(n14765), .ip2(n15093), .op(n15094) );
  nand2_1 U16469 ( .ip1(n21250), .ip2(n15094), .op(n15095) );
  nand2_1 U16470 ( .ip1(n15095), .ip2(\pipeline/md_resp_result [12]), .op(
        n15108) );
  nand2_1 U16471 ( .ip1(\pipeline/md/counter [3]), .ip2(
        \pipeline/md/counter [2]), .op(n18837) );
  nor2_1 U16472 ( .ip1(n21515), .ip2(n18837), .op(n18174) );
  nand2_1 U16473 ( .ip1(n21977), .ip2(n18174), .op(n15107) );
  inv_1 U16474 ( .ip(n15096), .op(n18072) );
  nor2_1 U16475 ( .ip1(\pipeline/md/result [43]), .ip2(n18072), .op(n18071) );
  inv_1 U16476 ( .ip(n18071), .op(n15098) );
  inv_1 U16477 ( .ip(\pipeline/md/result [44]), .op(n22588) );
  nand2_1 U16478 ( .ip1(n18071), .ip2(n22588), .op(n18163) );
  inv_1 U16479 ( .ip(n18163), .op(n15097) );
  not_ab_or_c_or_d U16480 ( .ip1(\pipeline/md/result [44]), .ip2(n15098), 
        .ip3(n15097), .ip4(n21505), .op(n15104) );
  nand2_1 U16481 ( .ip1(\pipeline/md/negate_output ), .ip2(n15099), .op(n15101) );
  nor2_1 U16482 ( .ip1(n15102), .ip2(n15101), .op(n15100) );
  not_ab_or_c_or_d U16483 ( .ip1(n15102), .ip2(n15101), .ip3(n21960), .ip4(
        n15100), .op(n15103) );
  not_ab_or_c_or_d U16484 ( .ip1(\pipeline/md/result [44]), .ip2(n21509), 
        .ip3(n15104), .ip4(n15103), .op(n15105) );
  or2_1 U16485 ( .ip1(n15105), .ip2(n21967), .op(n15106) );
  nand4_1 U16486 ( .ip1(n15109), .ip2(n15108), .ip3(n15107), .ip4(n15106), 
        .op(n8622) );
  or2_1 U16487 ( .ip1(n15111), .ip2(n15110), .op(n15113) );
  nand2_1 U16488 ( .ip1(n15113), .ip2(n15112), .op(n15114) );
  nor2_1 U16489 ( .ip1(\pipeline/md/b [13]), .ip2(n15114), .op(n15139) );
  or3_1 U16490 ( .ip1(n15139), .ip2(n15115), .ip3(n15116), .op(n15118) );
  nor2_1 U16491 ( .ip1(\pipeline/md_resp_result [13]), .ip2(n15118), .op(
        n15117) );
  nand2_1 U16492 ( .ip1(n21251), .ip2(n15117), .op(n15136) );
  nand2_1 U16493 ( .ip1(n20310), .ip2(n15118), .op(n15119) );
  nand2_1 U16494 ( .ip1(n21250), .ip2(n15119), .op(n15120) );
  nand2_1 U16495 ( .ip1(n15120), .ip2(\pipeline/md_resp_result [13]), .op(
        n15135) );
  nand2_1 U16496 ( .ip1(n20680), .ip2(n18174), .op(n15134) );
  or2_1 U16497 ( .ip1(n15121), .ip2(n21659), .op(n18159) );
  nor2_1 U16498 ( .ip1(n18157), .ip2(n18159), .op(n15125) );
  nor2_1 U16499 ( .ip1(n21960), .ip2(n21659), .op(n18081) );
  inv_1 U16500 ( .ip(n18081), .op(n21957) );
  nor2_1 U16501 ( .ip1(n15121), .ip2(n21957), .op(n15123) );
  nor2_1 U16502 ( .ip1(n21960), .ip2(n18157), .op(n15122) );
  nor2_1 U16503 ( .ip1(n15123), .ip2(n15122), .op(n15124) );
  nor2_1 U16504 ( .ip1(n15125), .ip2(n15124), .op(n15132) );
  nand2_1 U16505 ( .ip1(\pipeline/md/negate_output ), .ip2(n18163), .op(n15126) );
  nor2_1 U16506 ( .ip1(\pipeline/md/result [45]), .ip2(n15126), .op(n15128) );
  and2_1 U16507 ( .ip1(\pipeline/md/result [45]), .ip2(n15126), .op(n15127) );
  nor2_1 U16508 ( .ip1(n15128), .ip2(n15127), .op(n15129) );
  nor2_1 U16509 ( .ip1(n15129), .ip2(n21967), .op(n15130) );
  nor2_1 U16510 ( .ip1(n21972), .ip2(n15130), .op(n15131) );
  or2_1 U16511 ( .ip1(n15132), .ip2(n15131), .op(n15133) );
  nand4_1 U16512 ( .ip1(n15136), .ip2(n15135), .ip3(n15134), .ip4(n15133), 
        .op(n8621) );
  nor2_1 U16513 ( .ip1(\pipeline/md_resp_result [13]), .ip2(n15115), .op(
        n15138) );
  nor2_1 U16514 ( .ip1(n15138), .ip2(n15139), .op(n15137) );
  nor2_1 U16515 ( .ip1(\pipeline/md/b [14]), .ip2(n15137), .op(n18171) );
  inv_1 U16516 ( .ip(n18171), .op(n18175) );
  inv_1 U16517 ( .ip(n15138), .op(n15141) );
  inv_1 U16518 ( .ip(n15139), .op(n15140) );
  nand3_1 U16519 ( .ip1(\pipeline/md/b [14]), .ip2(n15141), .ip3(n15140), .op(
        n18176) );
  nand2_1 U16520 ( .ip1(n15142), .ip2(n18176), .op(n18170) );
  nand3_1 U16521 ( .ip1(\pipeline/md/b [15]), .ip2(n18175), .ip3(n18170), .op(
        n15148) );
  nand2_1 U16522 ( .ip1(n18175), .ip2(n18170), .op(n15143) );
  nand2_1 U16523 ( .ip1(n15144), .ip2(n15143), .op(n15164) );
  nand2_1 U16524 ( .ip1(n15148), .ip2(n15164), .op(n15145) );
  nand2_1 U16525 ( .ip1(n20310), .ip2(n15145), .op(n15146) );
  nand2_1 U16526 ( .ip1(n22738), .ip2(n15146), .op(n15147) );
  nand2_1 U16527 ( .ip1(\pipeline/md_resp_result [15]), .ip2(n15147), .op(
        n15162) );
  inv_1 U16528 ( .ip(n15148), .op(n15149) );
  nor2_1 U16529 ( .ip1(\pipeline/md_resp_result [15]), .ip2(n15149), .op(
        n15167) );
  nand3_1 U16530 ( .ip1(n22750), .ip2(n15167), .ip3(n15164), .op(n15161) );
  nand2_1 U16531 ( .ip1(\pipeline/md/negate_output ), .ip2(n15150), .op(n15152) );
  nor2_1 U16532 ( .ip1(n15153), .ip2(n15152), .op(n15151) );
  not_ab_or_c_or_d U16533 ( .ip1(n15153), .ip2(n15152), .ip3(n21960), .ip4(
        n15151), .op(n15158) );
  nor3_1 U16534 ( .ip1(\pipeline/md/result [46]), .ip2(
        \pipeline/md/result [45]), .ip3(n18163), .op(n15179) );
  nor3_1 U16535 ( .ip1(\pipeline/md/result [47]), .ip2(n15179), .ip3(n21966), 
        .op(n15156) );
  inv_1 U16536 ( .ip(n15179), .op(n15154) );
  inv_1 U16537 ( .ip(\pipeline/md/result [47]), .op(n22618) );
  not_ab_or_c_or_d U16538 ( .ip1(\pipeline/md/negate_output ), .ip2(n15154), 
        .ip3(n22618), .ip4(n21967), .op(n15155) );
  nor3_1 U16539 ( .ip1(n21972), .ip2(n15156), .ip3(n15155), .op(n15157) );
  or2_1 U16540 ( .ip1(n15158), .ip2(n15157), .op(n15160) );
  nand2_1 U16541 ( .ip1(n21671), .ip2(n18174), .op(n15159) );
  nand4_1 U16542 ( .ip1(n15162), .ip2(n15161), .ip3(n15160), .ip4(n15159), 
        .op(n8619) );
  nand2_1 U16543 ( .ip1(n18216), .ip2(\pipeline/md/counter [4]), .op(n18838)
         );
  nor2_1 U16544 ( .ip1(n15163), .ip2(n18838), .op(n20553) );
  nand2_1 U16545 ( .ip1(n21272), .ip2(n20553), .op(n15187) );
  inv_1 U16546 ( .ip(n15164), .op(n15168) );
  nor2_1 U16547 ( .ip1(n15168), .ip2(n15167), .op(n15165) );
  nor2_1 U16548 ( .ip1(\pipeline/md/b [16]), .ip2(n15165), .op(n18196) );
  nor3_1 U16549 ( .ip1(n15168), .ip2(n15167), .ip3(n15166), .op(n18195) );
  nor2_1 U16550 ( .ip1(\pipeline/md_resp_result [16]), .ip2(n18195), .op(
        n15169) );
  or2_1 U16551 ( .ip1(n18196), .ip2(n15169), .op(n15170) );
  nand2_1 U16552 ( .ip1(n15170), .ip2(n20010), .op(n15192) );
  inv_1 U16553 ( .ip(n15170), .op(n15171) );
  nand2_1 U16554 ( .ip1(\pipeline/md/b [17]), .ip2(n15171), .op(n15189) );
  nand2_1 U16555 ( .ip1(n15192), .ip2(n15189), .op(n15172) );
  nand2_1 U16556 ( .ip1(n20310), .ip2(n15172), .op(n15173) );
  nand2_1 U16557 ( .ip1(n22738), .ip2(n15173), .op(n15174) );
  nand2_1 U16558 ( .ip1(\pipeline/md_resp_result [17]), .ip2(n15174), .op(
        n15186) );
  inv_1 U16559 ( .ip(\pipeline/md_resp_result [17]), .op(n15190) );
  nand4_1 U16560 ( .ip1(n22750), .ip2(n15190), .ip3(n15192), .ip4(n15189), 
        .op(n15185) );
  nand2_1 U16561 ( .ip1(\pipeline/md/negate_output ), .ip2(n15175), .op(n15177) );
  nor2_1 U16562 ( .ip1(n15178), .ip2(n15177), .op(n15176) );
  not_ab_or_c_or_d U16563 ( .ip1(n15178), .ip2(n15177), .ip3(n21960), .ip4(
        n15176), .op(n15183) );
  inv_1 U16564 ( .ip(\pipeline/md/result [49]), .op(n22638) );
  nand2_1 U16565 ( .ip1(n15179), .ip2(n22618), .op(n18187) );
  nor2_1 U16566 ( .ip1(\pipeline/md/result [48]), .ip2(n18187), .op(n15201) );
  or2_1 U16567 ( .ip1(n15201), .ip2(n21659), .op(n18186) );
  nor2_1 U16568 ( .ip1(n22638), .ip2(n18186), .op(n15180) );
  not_ab_or_c_or_d U16569 ( .ip1(n22638), .ip2(n18186), .ip3(n15180), .ip4(
        n21967), .op(n15181) );
  nor2_1 U16570 ( .ip1(n21972), .ip2(n15181), .op(n15182) );
  or2_1 U16571 ( .ip1(n15183), .ip2(n15182), .op(n15184) );
  nand4_1 U16572 ( .ip1(n15187), .ip2(n15186), .ip3(n15185), .ip4(n15184), 
        .op(n8617) );
  nand2_1 U16573 ( .ip1(n15188), .ip2(n20553), .op(n15215) );
  nand2_1 U16574 ( .ip1(n15190), .ip2(n15189), .op(n15191) );
  nand2_1 U16575 ( .ip1(n15192), .ip2(n15191), .op(n15195) );
  inv_1 U16576 ( .ip(n15195), .op(n15193) );
  nor2_1 U16577 ( .ip1(\pipeline/md/b [18]), .ip2(n15193), .op(n15228) );
  nor2_1 U16578 ( .ip1(n15195), .ip2(n15194), .op(n15210) );
  or2_1 U16579 ( .ip1(n15228), .ip2(n15210), .op(n15196) );
  nand2_1 U16580 ( .ip1(n20310), .ip2(n15196), .op(n15197) );
  nand2_1 U16581 ( .ip1(n22738), .ip2(n15197), .op(n15198) );
  nand2_1 U16582 ( .ip1(\pipeline/md_resp_result [18]), .ip2(n15198), .op(
        n15214) );
  nor2_1 U16583 ( .ip1(n15199), .ip2(n21957), .op(n20546) );
  nor2_1 U16584 ( .ip1(n21960), .ip2(n20546), .op(n15206) );
  inv_1 U16585 ( .ip(\pipeline/md/result [50]), .op(n22651) );
  nor2_1 U16586 ( .ip1(n15200), .ip2(n22651), .op(n15204) );
  nand2_1 U16587 ( .ip1(n15201), .ip2(n22638), .op(n15202) );
  nor2_1 U16588 ( .ip1(\pipeline/md/result [50]), .ip2(n15202), .op(n20538) );
  not_ab_or_c_or_d U16589 ( .ip1(\pipeline/md/result [50]), .ip2(n15202), 
        .ip3(n20538), .ip4(n21505), .op(n15203) );
  not_ab_or_c_or_d U16590 ( .ip1(n15206), .ip2(n15205), .ip3(n15204), .ip4(
        n15203), .op(n15208) );
  nand2_1 U16591 ( .ip1(n20543), .ip2(n20546), .op(n15207) );
  nand2_1 U16592 ( .ip1(n15208), .ip2(n15207), .op(n15209) );
  nand2_1 U16593 ( .ip1(n20552), .ip2(n15209), .op(n15213) );
  nor2_1 U16594 ( .ip1(\pipeline/md_resp_result [18]), .ip2(n15210), .op(
        n15229) );
  inv_1 U16595 ( .ip(n15228), .op(n15211) );
  nand3_1 U16596 ( .ip1(n15229), .ip2(n22750), .ip3(n15211), .op(n15212) );
  nand4_1 U16597 ( .ip1(n15215), .ip2(n15214), .ip3(n15213), .ip4(n15212), 
        .op(n8616) );
  inv_1 U16598 ( .ip(\pipeline/md/result [51]), .op(n15216) );
  nand2_1 U16599 ( .ip1(n20538), .ip2(n15216), .op(n18256) );
  nor2_1 U16600 ( .ip1(\pipeline/md/result [52]), .ip2(n18256), .op(n20453) );
  inv_1 U16601 ( .ip(\pipeline/md/result [53]), .op(n22679) );
  nand2_1 U16602 ( .ip1(n20453), .ip2(n22679), .op(n18100) );
  nor2_1 U16603 ( .ip1(\pipeline/md/result [54]), .ip2(n18100), .op(n18117) );
  inv_1 U16604 ( .ip(\pipeline/md/result [55]), .op(n22700) );
  nand2_1 U16605 ( .ip1(n18117), .ip2(n22700), .op(n21969) );
  or2_1 U16606 ( .ip1(\pipeline/md/result [56]), .ip2(n21969), .op(n15217) );
  nor2_1 U16607 ( .ip1(n15217), .ip2(\pipeline/md/result [57]), .op(n15260) );
  not_ab_or_c_or_d U16608 ( .ip1(\pipeline/md/result [57]), .ip2(n15217), 
        .ip3(n15260), .ip4(n21505), .op(n15225) );
  inv_1 U16609 ( .ip(n21958), .op(n21955) );
  nor2_1 U16610 ( .ip1(n21955), .ip2(n21959), .op(n15218) );
  nor2_1 U16611 ( .ip1(n15218), .ip2(n21659), .op(n15219) );
  xor2_1 U16612 ( .ip1(n15220), .ip2(n15219), .op(n15221) );
  nor2_1 U16613 ( .ip1(n15221), .ip2(n15265), .op(n15224) );
  inv_1 U16614 ( .ip(\pipeline/md/result [57]), .op(n15222) );
  nor2_1 U16615 ( .ip1(n15267), .ip2(n15222), .op(n15223) );
  not_ab_or_c_or_d U16616 ( .ip1(n20552), .ip2(n15225), .ip3(n15224), .ip4(
        n15223), .op(n15259) );
  inv_1 U16617 ( .ip(\pipeline/md_resp_result [22]), .op(n15237) );
  nor2_1 U16618 ( .ip1(n15229), .ip2(n15228), .op(n15226) );
  nor2_1 U16619 ( .ip1(\pipeline/md/b [19]), .ip2(n15226), .op(n20556) );
  nor3_1 U16620 ( .ip1(n15229), .ip2(n15228), .ip3(n15227), .op(n20555) );
  nor2_1 U16621 ( .ip1(\pipeline/md_resp_result [19]), .ip2(n20555), .op(
        n15230) );
  nor2_1 U16622 ( .ip1(n20556), .ip2(n15230), .op(n15231) );
  nor2_1 U16623 ( .ip1(\pipeline/md/b [20]), .ip2(n15231), .op(n18264) );
  inv_1 U16624 ( .ip(n15231), .op(n15232) );
  nor2_1 U16625 ( .ip1(n20577), .ip2(n15232), .op(n18263) );
  nor2_1 U16626 ( .ip1(\pipeline/md_resp_result [20]), .ip2(n18263), .op(
        n15233) );
  nor2_1 U16627 ( .ip1(n18264), .ip2(n15233), .op(n15234) );
  nor2_1 U16628 ( .ip1(\pipeline/md/b [21]), .ip2(n15234), .op(n20463) );
  inv_1 U16629 ( .ip(n15234), .op(n15235) );
  nor2_1 U16630 ( .ip1(n20590), .ip2(n15235), .op(n20462) );
  nor2_1 U16631 ( .ip1(\pipeline/md_resp_result [21]), .ip2(n20462), .op(
        n15236) );
  nor2_1 U16632 ( .ip1(n20463), .ip2(n15236), .op(n15238) );
  nor2_1 U16633 ( .ip1(\pipeline/md/b [22]), .ip2(n15238), .op(n18109) );
  or2_1 U16634 ( .ip1(n15237), .ip2(n18109), .op(n15239) );
  nand2_1 U16635 ( .ip1(\pipeline/md/b [22]), .ip2(n15238), .op(n18110) );
  nand2_1 U16636 ( .ip1(n15239), .ip2(n18110), .op(n15240) );
  nor2_1 U16637 ( .ip1(\pipeline/md/b [23]), .ip2(n15240), .op(n18132) );
  inv_1 U16638 ( .ip(n15240), .op(n15241) );
  nor2_1 U16639 ( .ip1(n15242), .ip2(n15241), .op(n18131) );
  nor2_1 U16640 ( .ip1(\pipeline/md_resp_result [23]), .ip2(n18131), .op(
        n15243) );
  nor2_1 U16641 ( .ip1(n18132), .ip2(n15243), .op(n15244) );
  nor2_1 U16642 ( .ip1(\pipeline/md/b [24]), .ip2(n15244), .op(n21979) );
  nor2_1 U16643 ( .ip1(\pipeline/md_resp_result [24]), .ip2(n15245), .op(
        n15246) );
  nor2_1 U16644 ( .ip1(n21979), .ip2(n15246), .op(n15247) );
  nand2_1 U16645 ( .ip1(\pipeline/md/b [25]), .ip2(n15247), .op(n15253) );
  inv_1 U16646 ( .ip(n15247), .op(n15248) );
  nand2_1 U16647 ( .ip1(n15249), .ip2(n15248), .op(n15271) );
  nand2_1 U16648 ( .ip1(n15253), .ip2(n15271), .op(n15250) );
  nand2_1 U16649 ( .ip1(n20310), .ip2(n15250), .op(n15251) );
  nand2_1 U16650 ( .ip1(n22738), .ip2(n15251), .op(n15252) );
  nand2_1 U16651 ( .ip1(\pipeline/md_resp_result [25]), .ip2(n15252), .op(
        n15258) );
  inv_1 U16652 ( .ip(n22750), .op(n22755) );
  inv_1 U16653 ( .ip(n15253), .op(n15254) );
  nor2_1 U16654 ( .ip1(\pipeline/md_resp_result [25]), .ip2(n15254), .op(
        n15274) );
  nand3_1 U16655 ( .ip1(n22750), .ip2(n15274), .ip3(n15271), .op(n15257) );
  nor2_1 U16656 ( .ip1(n15255), .ip2(n18838), .op(n21978) );
  nand2_1 U16657 ( .ip1(n21978), .ip2(n20680), .op(n15256) );
  nand4_1 U16658 ( .ip1(n15259), .ip2(n15258), .ip3(n15257), .ip4(n15256), 
        .op(n8609) );
  inv_1 U16659 ( .ip(n15260), .op(n20296) );
  or2_1 U16660 ( .ip1(\pipeline/md/result [58]), .ip2(n20296), .op(n15261) );
  nor2_1 U16661 ( .ip1(n15261), .ip2(\pipeline/md/result [59]), .op(n19017) );
  not_ab_or_c_or_d U16662 ( .ip1(\pipeline/md/result [59]), .ip2(n15261), 
        .ip3(n19017), .ip4(n21505), .op(n15270) );
  nor2_1 U16663 ( .ip1(n15262), .ip2(n21659), .op(n15263) );
  xor2_1 U16664 ( .ip1(n15264), .ip2(n15263), .op(n15266) );
  nor2_1 U16665 ( .ip1(n15266), .ip2(n15265), .op(n15269) );
  inv_1 U16666 ( .ip(\pipeline/md/result [59]), .op(n22722) );
  nor2_1 U16667 ( .ip1(n15267), .ip2(n22722), .op(n15268) );
  not_ab_or_c_or_d U16668 ( .ip1(n20552), .ip2(n15270), .ip3(n15269), .ip4(
        n15268), .op(n15286) );
  inv_1 U16669 ( .ip(n15271), .op(n15275) );
  nor2_1 U16670 ( .ip1(n15275), .ip2(n15274), .op(n15272) );
  nor2_1 U16671 ( .ip1(\pipeline/md/b [26]), .ip2(n15272), .op(n20308) );
  nor3_1 U16672 ( .ip1(n15275), .ip2(n15274), .ip3(n15273), .op(n20307) );
  nor2_1 U16673 ( .ip1(\pipeline/md_resp_result [26]), .ip2(n20307), .op(
        n15276) );
  nor2_1 U16674 ( .ip1(n20308), .ip2(n15276), .op(n15277) );
  nor2_1 U16675 ( .ip1(\pipeline/md/b [27]), .ip2(n15277), .op(n18841) );
  inv_1 U16676 ( .ip(n15277), .op(n15278) );
  nor2_1 U16677 ( .ip1(n15279), .ip2(n15278), .op(n18839) );
  or2_1 U16678 ( .ip1(n18841), .ip2(n18839), .op(n15280) );
  nand2_1 U16679 ( .ip1(n20310), .ip2(n15280), .op(n15281) );
  nand2_1 U16680 ( .ip1(n22738), .ip2(n15281), .op(n15282) );
  nand2_1 U16681 ( .ip1(\pipeline/md_resp_result [27]), .ip2(n15282), .op(
        n15285) );
  or4_1 U16682 ( .ip1(\pipeline/md_resp_result [27]), .ip2(n18841), .ip3(
        n18839), .ip4(n22755), .op(n15284) );
  nand2_1 U16683 ( .ip1(n21671), .ip2(n21978), .op(n15283) );
  nand4_1 U16684 ( .ip1(n15286), .ip2(n15285), .ip3(n15284), .ip4(n15283), 
        .op(n8607) );
  nand2_1 U16685 ( .ip1(n21683), .ip2(n22665), .op(n21680) );
  nand2_1 U16686 ( .ip1(n17747), .ip2(n21680), .op(n15288) );
  nand2_1 U16687 ( .ip1(\pipeline/md/counter [1]), .ip2(n22665), .op(n15287)
         );
  nand4_1 U16688 ( .ip1(n21683), .ip2(n15289), .ip3(n15288), .ip4(n15287), 
        .op(n8537) );
  mux2_1 U16689 ( .ip1(n15291), .ip2(n15290), .s(n17399), .op(n17298) );
  mux2_1 U16690 ( .ip1(\pipeline/dmem_type[2] ), .ip2(n16478), .s(
        dmem_hsize[0]), .op(n21686) );
  nand2_1 U16691 ( .ip1(n22069), .ip2(n21686), .op(n21414) );
  nor2_1 U16692 ( .ip1(n21414), .ip2(n21683), .op(n21360) );
  nor2_1 U16693 ( .ip1(n22053), .ip2(n22055), .op(n17299) );
  inv_1 U16694 ( .ip(n17299), .op(n15292) );
  nand3_1 U16695 ( .ip1(n17298), .ip2(n21360), .ip3(n15292), .op(n15298) );
  nand2_1 U16696 ( .ip1(n21440), .ip2(\pipeline/md/b [34]), .op(n15297) );
  inv_1 U16697 ( .ip(n17298), .op(n22057) );
  inv_1 U16698 ( .ip(n21414), .op(n21427) );
  nor2_1 U16699 ( .ip1(n21427), .ip2(n21683), .op(n21400) );
  inv_1 U16700 ( .ip(n21400), .op(n21409) );
  inv_1 U16701 ( .ip(n21683), .op(n22042) );
  nand2_1 U16702 ( .ip1(n22042), .ip2(n17299), .op(n15293) );
  nand2_1 U16703 ( .ip1(n21409), .ip2(n15293), .op(n15294) );
  nand2_1 U16704 ( .ip1(n22057), .ip2(n15294), .op(n15296) );
  inv_1 U16705 ( .ip(n21680), .op(n21496) );
  buf_1 U16706 ( .ip(n21496), .op(n21493) );
  nand2_1 U16707 ( .ip1(n21493), .ip2(\pipeline/md/b [33]), .op(n15295) );
  nand4_1 U16708 ( .ip1(n15298), .ip2(n15297), .ip3(n15296), .ip4(n15295), 
        .op(n8368) );
  nand2_1 U16709 ( .ip1(n21493), .ip2(\pipeline/md/b [32]), .op(n15306) );
  nand2_1 U16710 ( .ip1(n21440), .ip2(\pipeline/md/b [33]), .op(n15305) );
  inv_1 U16711 ( .ip(n22055), .op(n15299) );
  nand3_1 U16712 ( .ip1(n15299), .ip2(n21360), .ip3(n22053), .op(n15304) );
  inv_1 U16713 ( .ip(n22053), .op(n15300) );
  nand2_1 U16714 ( .ip1(n15300), .ip2(n22042), .op(n15301) );
  nand2_1 U16715 ( .ip1(n21409), .ip2(n15301), .op(n15302) );
  nand2_1 U16716 ( .ip1(n22055), .ip2(n15302), .op(n15303) );
  nand4_1 U16717 ( .ip1(n15306), .ip2(n15305), .ip3(n15304), .ip4(n15303), 
        .op(n8367) );
  inv_1 U16718 ( .ip(htif_pcr_resp_valid), .op(htif_pcr_req_ready) );
  nand2_1 U16719 ( .ip1(htif_pcr_req_valid), .ip2(htif_pcr_req_ready), .op(
        n22476) );
  inv_1 U16720 ( .ip(n22476), .op(n15307) );
  nand2_1 U16721 ( .ip1(n15307), .ip2(htif_pcr_req_rw), .op(n15725) );
  inv_1 U16722 ( .ip(n15725), .op(n16369) );
  or2_1 U16723 ( .ip1(\pipeline/csr/system_wen ), .ip2(n16369), .op(n20965) );
  nor3_1 U16724 ( .ip1(\pipeline/inst_DX [27]), .ip2(n22120), .ip3(n22121), 
        .op(n22104) );
  nand3_1 U16725 ( .ip1(n22104), .ip2(n15324), .ip3(n15308), .op(n15331) );
  nor2_1 U16726 ( .ip1(\pipeline/inst_DX [25]), .ip2(n15331), .op(n22098) );
  nand2_1 U16727 ( .ip1(\pipeline/inst_DX [26]), .ip2(n22098), .op(n22110) );
  nor2_1 U16728 ( .ip1(n15309), .ip2(n22110), .op(n16396) );
  nand2_1 U16729 ( .ip1(n20965), .ip2(n16396), .op(n15857) );
  inv_1 U16730 ( .ip(n15857), .op(n16410) );
  inv_1 U16731 ( .ip(n15310), .op(n17884) );
  nand2_1 U16732 ( .ip1(n17884), .ip2(n17786), .op(n17782) );
  nor2_1 U16733 ( .ip1(n17782), .ip2(n17819), .op(n22091) );
  inv_1 U16734 ( .ip(n15311), .op(n15353) );
  nor2_1 U16735 ( .ip1(n15353), .ip2(n15312), .op(n15313) );
  and2_1 U16736 ( .ip1(n22091), .ip2(n15313), .op(n22896) );
  nand2_1 U16737 ( .ip1(n22896), .ip2(dmem_hsize[1]), .op(n15314) );
  and2_1 U16738 ( .ip1(\pipeline/csr/system_wen ), .ip2(n15725), .op(n15355)
         );
  nand2_1 U16739 ( .ip1(n15314), .ip2(n15355), .op(n16019) );
  nand2_1 U16740 ( .ip1(n16019), .ip2(n20965), .op(n17949) );
  and2_1 U16741 ( .ip1(n17949), .ip2(n17765), .op(n16368) );
  nand2_1 U16742 ( .ip1(n16368), .ip2(n15356), .op(n15362) );
  and2_1 U16743 ( .ip1(n16369), .ip2(htif_pcr_req_data[20]), .op(n15360) );
  inv_1 U16744 ( .ip(n22119), .op(n15674) );
  nor2_1 U16745 ( .ip1(n15674), .ip2(n22110), .op(n17828) );
  inv_1 U16746 ( .ip(n15315), .op(n17630) );
  nand2_1 U16747 ( .ip1(\pipeline/inst_DX [30]), .ip2(n15324), .op(n15321) );
  nor2_1 U16748 ( .ip1(\pipeline/inst_DX [25]), .ip2(n15321), .op(n22103) );
  nand3_1 U16749 ( .ip1(n17630), .ip2(n22103), .ip3(n22104), .op(n18439) );
  inv_1 U16750 ( .ip(n18439), .op(n15316) );
  nand2_1 U16751 ( .ip1(\pipeline/inst_DX [26]), .ip2(n15316), .op(n18440) );
  nor2_1 U16752 ( .ip1(n15340), .ip2(n18440), .op(n16310) );
  inv_1 U16753 ( .ip(n16310), .op(n16338) );
  inv_1 U16754 ( .ip(\pipeline/csr/mtime_full [52]), .op(n22196) );
  nor2_1 U16755 ( .ip1(n16338), .ip2(n22196), .op(n15320) );
  nand2_1 U16756 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [20]), .op(n15318) );
  inv_1 U16757 ( .ip(n22109), .op(n15731) );
  nor2_1 U16758 ( .ip1(n15731), .ip2(n22110), .op(n17305) );
  nand2_1 U16759 ( .ip1(\pipeline/epc [20]), .ip2(n17305), .op(n15317) );
  nand2_1 U16760 ( .ip1(n15318), .ip2(n15317), .op(n15319) );
  not_ab_or_c_or_d U16761 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [20]), 
        .ip3(n15320), .ip4(n15319), .op(n15351) );
  inv_1 U16762 ( .ip(n15330), .op(n15325) );
  nor2_1 U16763 ( .ip1(n15325), .ip2(n15321), .op(n15322) );
  nand4_1 U16764 ( .ip1(\pipeline/inst_DX [28]), .ip2(\pipeline/inst_DX [29]), 
        .ip3(\pipeline/inst_DX [27]), .ip4(n15322), .op(n22099) );
  or2_1 U16765 ( .ip1(n15674), .ip2(n22099), .op(n17843) );
  inv_1 U16766 ( .ip(n17843), .op(n22096) );
  xor2_1 U16767 ( .ip1(\pipeline/inst_DX [30]), .ip2(n22120), .op(n15323) );
  nor4_1 U16768 ( .ip1(\pipeline/inst_DX [29]), .ip2(n15325), .ip3(n15324), 
        .ip4(n15323), .op(n22092) );
  nand3_1 U16769 ( .ip1(n15338), .ip2(n22092), .ip3(n15339), .op(n16380) );
  inv_1 U16770 ( .ip(\pipeline/csr/instret_full [20]), .op(n19541) );
  nor2_1 U16771 ( .ip1(n16380), .ip2(n19541), .op(n15328) );
  nor2_1 U16772 ( .ip1(n15731), .ip2(n22099), .op(n16383) );
  nand4_1 U16773 ( .ip1(n15330), .ip2(\pipeline/imm[31] ), .ip3(
        \pipeline/inst_DX [30]), .ip4(n22104), .op(n22100) );
  nor2_1 U16774 ( .ip1(n15674), .ip2(n22100), .op(n15434) );
  nor3_1 U16775 ( .ip1(\pipeline/inst_DX [26]), .ip2(n15340), .ip3(n18439), 
        .op(n16382) );
  inv_1 U16776 ( .ip(n16382), .op(n15971) );
  inv_1 U16777 ( .ip(\pipeline/csr/mtime_full [20]), .op(n19658) );
  nor2_1 U16778 ( .ip1(n15971), .ip2(n19658), .op(n15326) );
  ab_or_c_or_d U16779 ( .ip1(n16383), .ip2(\pipeline/csr/from_host [20]), 
        .ip3(n15434), .ip4(n15326), .op(n15327) );
  not_ab_or_c_or_d U16780 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [20]), 
        .ip3(n15328), .ip4(n15327), .op(n15350) );
  inv_1 U16781 ( .ip(n22097), .op(n15347) );
  inv_1 U16782 ( .ip(n15331), .op(n15329) );
  nand2_1 U16783 ( .ip1(n15330), .ip2(n15329), .op(n15673) );
  nor2_1 U16784 ( .ip1(n15347), .ip2(n15673), .op(n18144) );
  nand2_1 U16785 ( .ip1(\pipeline/csr/mie [20]), .ip2(n18144), .op(n15336) );
  or2_1 U16786 ( .ip1(n15332), .ip2(n15331), .op(n22105) );
  or2_1 U16787 ( .ip1(n15731), .ip2(n22105), .op(n15533) );
  inv_1 U16788 ( .ip(n15533), .op(n17812) );
  nand2_1 U16789 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [20]), .op(n15335) );
  nand2_1 U16790 ( .ip1(\pipeline/inst_DX [27]), .ip2(n22092), .op(n17628) );
  nor2_1 U16791 ( .ip1(n15674), .ip2(n17628), .op(n16387) );
  nand2_1 U16792 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [52]), .op(
        n15334) );
  nor2_1 U16793 ( .ip1(n15731), .ip2(n15673), .op(n17364) );
  nand2_1 U16794 ( .ip1(\pipeline/csr/mtvec [20]), .ip2(n17364), .op(n15333)
         );
  nand4_1 U16795 ( .ip1(n15336), .ip2(n15335), .ip3(n15334), .ip4(n15333), 
        .op(n15346) );
  inv_1 U16796 ( .ip(n22094), .op(n15337) );
  nand3_1 U16797 ( .ip1(n15337), .ip2(n22092), .ip3(n15339), .op(n18456) );
  nor2_1 U16798 ( .ip1(n15340), .ip2(n18456), .op(n16370) );
  nand2_1 U16799 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [20]), .op(
        n15344) );
  inv_1 U16800 ( .ip(n15338), .op(n22093) );
  nor2_1 U16801 ( .ip1(n22093), .ip2(n17628), .op(n16371) );
  nand2_1 U16802 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [52]), .op(
        n15343) );
  nand3_1 U16803 ( .ip1(n17630), .ip2(n22092), .ip3(n15339), .op(n17597) );
  or2_1 U16804 ( .ip1(n15340), .ip2(n17597), .op(n15538) );
  inv_1 U16805 ( .ip(n15538), .op(n16372) );
  nand2_1 U16806 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [20]), .op(
        n15342) );
  nor2_1 U16807 ( .ip1(n15731), .ip2(n17628), .op(n16373) );
  nand2_1 U16808 ( .ip1(n16373), .ip2(\pipeline/csr/time_full [52]), .op(
        n15341) );
  nand4_1 U16809 ( .ip1(n15344), .ip2(n15343), .ip3(n15342), .ip4(n15341), 
        .op(n15345) );
  nor2_1 U16810 ( .ip1(n15346), .ip2(n15345), .op(n15349) );
  nor2_1 U16811 ( .ip1(n15347), .ip2(n22110), .op(n19599) );
  nand2_1 U16812 ( .ip1(ext_interrupts[12]), .ip2(n19599), .op(n15348) );
  and4_1 U16813 ( .ip1(n15351), .ip2(n15350), .ip3(n15349), .ip4(n15348), .op(
        n19555) );
  nor2_1 U16814 ( .ip1(n15353), .ip2(n15352), .op(n15354) );
  and2_1 U16815 ( .ip1(n22091), .ip2(n15354), .op(n22898) );
  nand2_1 U16816 ( .ip1(n22898), .ip2(n15355), .op(n16401) );
  nor2_1 U16817 ( .ip1(n15356), .ip2(n16401), .op(n15357) );
  nor2_1 U16818 ( .ip1(n17765), .ip2(n16401), .op(n16403) );
  nor2_1 U16819 ( .ip1(n15357), .ip2(n16403), .op(n15358) );
  nor2_1 U16820 ( .ip1(n19555), .ip2(n15358), .op(n15359) );
  nor2_1 U16821 ( .ip1(n15360), .ip2(n15359), .op(n15361) );
  nand2_1 U16822 ( .ip1(n15362), .ip2(n15361), .op(n19549) );
  nand2_1 U16823 ( .ip1(n16410), .ip2(n19549), .op(n15368) );
  nor2_1 U16824 ( .ip1(n16410), .ip2(n21082), .op(n16411) );
  nand2_1 U16825 ( .ip1(\pipeline/csr/mbadaddr [20]), .ip2(n16411), .op(n15367) );
  inv_1 U16826 ( .ip(\pipeline/ctrl/had_ex_WB ), .op(n16056) );
  nor4_1 U16827 ( .ip1(\pipeline/ctrl/prev_ex_code_WB [3]), .ip2(
        \pipeline/ctrl/prev_ex_code_WB [1]), .ip3(
        \pipeline/ctrl/prev_ex_code_WB [0]), .ip4(n16056), .op(n15363) );
  nor3_1 U16828 ( .ip1(n20972), .ip2(n16410), .ip3(n15363), .op(n16412) );
  nand2_1 U16829 ( .ip1(\pipeline/alu_out_WB [20]), .ip2(n16412), .op(n15366)
         );
  inv_1 U16830 ( .ip(n15363), .op(n15364) );
  nor2_1 U16831 ( .ip1(n16410), .ip2(n15364), .op(n16413) );
  nand2_1 U16832 ( .ip1(n16413), .ip2(\pipeline/PC_WB [20]), .op(n15365) );
  nand4_1 U16833 ( .ip1(n15368), .ip2(n15367), .ip3(n15366), .ip4(n15365), 
        .op(n8680) );
  nand2_1 U16834 ( .ip1(n16368), .ip2(n15369), .op(n15396) );
  nand2_1 U16835 ( .ip1(n16369), .ip2(htif_pcr_req_data[22]), .op(n15395) );
  inv_1 U16836 ( .ip(n16403), .op(n16337) );
  inv_1 U16837 ( .ip(n16401), .op(n16335) );
  nand2_1 U16838 ( .ip1(n16335), .ip2(n20599), .op(n15370) );
  nand2_1 U16839 ( .ip1(n16337), .ip2(n15370), .op(n15393) );
  nand2_1 U16840 ( .ip1(ext_interrupts[14]), .ip2(n19599), .op(n15392) );
  nand2_1 U16841 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [54]), .op(
        n15374) );
  inv_1 U16842 ( .ip(n16380), .op(n16301) );
  nand2_1 U16843 ( .ip1(n16301), .ip2(\pipeline/csr/instret_full [22]), .op(
        n15373) );
  nand2_1 U16844 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [22]), .op(n15372)
         );
  nand2_1 U16845 ( .ip1(n16383), .ip2(\pipeline/csr/from_host [22]), .op(
        n15371) );
  nand4_1 U16846 ( .ip1(n15374), .ip2(n15373), .ip3(n15372), .ip4(n15371), 
        .op(n15378) );
  nand2_1 U16847 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [22]), .op(n15376) );
  nand2_1 U16848 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [22]), .op(n15375) );
  nand2_1 U16849 ( .ip1(n15376), .ip2(n15375), .op(n15377) );
  not_ab_or_c_or_d U16850 ( .ip1(n16310), .ip2(\pipeline/csr/mtime_full [54]), 
        .ip3(n15378), .ip4(n15377), .op(n15391) );
  nand2_1 U16851 ( .ip1(\pipeline/csr/mie [22]), .ip2(n18144), .op(n15382) );
  nand2_1 U16852 ( .ip1(n16382), .ip2(\pipeline/csr/mtime_full [22]), .op(
        n15381) );
  nand2_1 U16853 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [22]), .op(n15380) );
  nand2_1 U16854 ( .ip1(\pipeline/csr/mtvec [22]), .ip2(n17364), .op(n15379)
         );
  nand4_1 U16855 ( .ip1(n15382), .ip2(n15381), .ip3(n15380), .ip4(n15379), 
        .op(n15388) );
  nand2_1 U16856 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [54]), .op(
        n15386) );
  nand2_1 U16857 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [22]), .op(
        n15385) );
  nand2_1 U16858 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [22]), .op(
        n15384) );
  nand2_1 U16859 ( .ip1(n16373), .ip2(\pipeline/csr/time_full [54]), .op(
        n15383) );
  nand4_1 U16860 ( .ip1(n15386), .ip2(n15385), .ip3(n15384), .ip4(n15383), 
        .op(n15387) );
  nor2_1 U16861 ( .ip1(n15388), .ip2(n15387), .op(n15390) );
  nand2_1 U16862 ( .ip1(\pipeline/epc [22]), .ip2(n17305), .op(n15389) );
  nand4_1 U16863 ( .ip1(n15392), .ip2(n15391), .ip3(n15390), .ip4(n15389), 
        .op(n20105) );
  nand2_1 U16864 ( .ip1(n15393), .ip2(n20105), .op(n15394) );
  nand3_1 U16865 ( .ip1(n15396), .ip2(n15395), .ip3(n15394), .op(n20100) );
  nand2_1 U16866 ( .ip1(n16410), .ip2(n20100), .op(n15400) );
  nand2_1 U16867 ( .ip1(\pipeline/csr/mbadaddr [22]), .ip2(n16411), .op(n15399) );
  nand2_1 U16868 ( .ip1(\pipeline/alu_out_WB [22]), .ip2(n16412), .op(n15398)
         );
  nand2_1 U16869 ( .ip1(n16413), .ip2(\pipeline/PC_WB [22]), .op(n15397) );
  nand4_1 U16870 ( .ip1(n15400), .ip2(n15399), .ip3(n15398), .ip4(n15397), 
        .op(n8678) );
  nand2_1 U16871 ( .ip1(n16368), .ip2(n15401), .op(n15428) );
  nand2_1 U16872 ( .ip1(n16369), .ip2(htif_pcr_req_data[23]), .op(n15427) );
  nand2_1 U16873 ( .ip1(n16335), .ip2(n20278), .op(n15402) );
  nand2_1 U16874 ( .ip1(n16337), .ip2(n15402), .op(n15425) );
  nand2_1 U16875 ( .ip1(ext_interrupts[15]), .ip2(n19599), .op(n15424) );
  nand2_1 U16876 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [55]), .op(
        n15406) );
  nand2_1 U16877 ( .ip1(n16301), .ip2(\pipeline/csr/instret_full [23]), .op(
        n15405) );
  nand2_1 U16878 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [23]), .op(n15404)
         );
  nand2_1 U16879 ( .ip1(n16383), .ip2(\pipeline/csr/from_host [23]), .op(
        n15403) );
  nand4_1 U16880 ( .ip1(n15406), .ip2(n15405), .ip3(n15404), .ip4(n15403), 
        .op(n15410) );
  nand2_1 U16881 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [23]), .op(n15408) );
  nand2_1 U16882 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [23]), .op(n15407) );
  nand2_1 U16883 ( .ip1(n15408), .ip2(n15407), .op(n15409) );
  not_ab_or_c_or_d U16884 ( .ip1(n16310), .ip2(\pipeline/csr/mtime_full [55]), 
        .ip3(n15410), .ip4(n15409), .op(n15423) );
  nand2_1 U16885 ( .ip1(\pipeline/csr/mie [23]), .ip2(n18144), .op(n15414) );
  nand2_1 U16886 ( .ip1(n16382), .ip2(\pipeline/csr/mtime_full [23]), .op(
        n15413) );
  nand2_1 U16887 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [23]), .op(n15412) );
  nand2_1 U16888 ( .ip1(\pipeline/csr/mtvec [23]), .ip2(n17364), .op(n15411)
         );
  nand4_1 U16889 ( .ip1(n15414), .ip2(n15413), .ip3(n15412), .ip4(n15411), 
        .op(n15420) );
  nand2_1 U16890 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [55]), .op(
        n15418) );
  nand2_1 U16891 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [23]), .op(
        n15417) );
  nand2_1 U16892 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [23]), .op(
        n15416) );
  nand2_1 U16893 ( .ip1(n16373), .ip2(\pipeline/csr/time_full [55]), .op(
        n15415) );
  nand4_1 U16894 ( .ip1(n15418), .ip2(n15417), .ip3(n15416), .ip4(n15415), 
        .op(n15419) );
  nor2_1 U16895 ( .ip1(n15420), .ip2(n15419), .op(n15422) );
  nand2_1 U16896 ( .ip1(\pipeline/epc [23]), .ip2(n17305), .op(n15421) );
  nand4_1 U16897 ( .ip1(n15424), .ip2(n15423), .ip3(n15422), .ip4(n15421), 
        .op(n20145) );
  nand2_1 U16898 ( .ip1(n15425), .ip2(n20145), .op(n15426) );
  nand3_1 U16899 ( .ip1(n15428), .ip2(n15427), .ip3(n15426), .op(n22274) );
  nand2_1 U16900 ( .ip1(n16410), .ip2(n22274), .op(n15432) );
  nand2_1 U16901 ( .ip1(\pipeline/csr/mbadaddr [23]), .ip2(n16411), .op(n15431) );
  nand2_1 U16902 ( .ip1(\pipeline/alu_out_WB [23]), .ip2(n16412), .op(n15430)
         );
  nand2_1 U16903 ( .ip1(n16413), .ip2(\pipeline/PC_WB [23]), .op(n15429) );
  nand4_1 U16904 ( .ip1(n15432), .ip2(n15431), .ip3(n15430), .ip4(n15429), 
        .op(n8677) );
  inv_1 U16905 ( .ip(n15433), .op(n19748) );
  nand2_1 U16906 ( .ip1(n16368), .ip2(n19748), .op(n15462) );
  and2_1 U16907 ( .ip1(n16369), .ip2(htif_pcr_req_data[8]), .op(n15460) );
  inv_1 U16908 ( .ip(\pipeline/csr/mtime_full [8]), .op(n19637) );
  nor2_1 U16909 ( .ip1(n15971), .ip2(n19637), .op(n15435) );
  not_ab_or_c_or_d U16910 ( .ip1(n16383), .ip2(\pipeline/csr/from_host [8]), 
        .ip3(n15435), .ip4(n15434), .op(n15438) );
  nand2_1 U16911 ( .ip1(n16301), .ip2(\pipeline/csr/instret_full [8]), .op(
        n15437) );
  nand2_1 U16912 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [8]), .op(n15436)
         );
  nand3_1 U16913 ( .ip1(n15438), .ip2(n15437), .ip3(n15436), .op(n15450) );
  nand2_1 U16914 ( .ip1(\pipeline/csr/mie [8]), .ip2(n18144), .op(n15442) );
  nand2_1 U16915 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [8]), .op(n15441)
         );
  nand2_1 U16916 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [40]), .op(
        n15440) );
  nand2_1 U16917 ( .ip1(\pipeline/csr/mtvec [8]), .ip2(n17364), .op(n15439) );
  nand4_1 U16918 ( .ip1(n15442), .ip2(n15441), .ip3(n15440), .ip4(n15439), 
        .op(n15448) );
  nand2_1 U16919 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [8]), .op(
        n15446) );
  nand2_1 U16920 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [40]), .op(
        n15445) );
  nand2_1 U16921 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [8]), .op(n15444) );
  nand2_1 U16922 ( .ip1(n16373), .ip2(\pipeline/csr/time_full [40]), .op(
        n15443) );
  nand4_1 U16923 ( .ip1(n15446), .ip2(n15445), .ip3(n15444), .ip4(n15443), 
        .op(n15447) );
  or2_1 U16924 ( .ip1(n15448), .ip2(n15447), .op(n15449) );
  not_ab_or_c_or_d U16925 ( .ip1(n19599), .ip2(ext_interrupts[0]), .ip3(n15450), .ip4(n15449), .op(n15456) );
  inv_1 U16926 ( .ip(\pipeline/csr/mtime_full [40]), .op(n18450) );
  nor2_1 U16927 ( .ip1(n16338), .ip2(n18450), .op(n15454) );
  nand2_1 U16928 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [8]), .op(n15452)
         );
  nand2_1 U16929 ( .ip1(\pipeline/epc [8]), .ip2(n17305), .op(n15451) );
  nand2_1 U16930 ( .ip1(n15452), .ip2(n15451), .op(n15453) );
  not_ab_or_c_or_d U16931 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [8]), 
        .ip3(n15454), .ip4(n15453), .op(n15455) );
  and2_1 U16932 ( .ip1(n15456), .ip2(n15455), .op(n19745) );
  nor2_1 U16933 ( .ip1(n19748), .ip2(n16401), .op(n15457) );
  nor2_1 U16934 ( .ip1(n15457), .ip2(n16403), .op(n15458) );
  nor2_1 U16935 ( .ip1(n19745), .ip2(n15458), .op(n15459) );
  nor2_1 U16936 ( .ip1(n15460), .ip2(n15459), .op(n15461) );
  and2_1 U16937 ( .ip1(n15462), .ip2(n15461), .op(n19700) );
  inv_1 U16938 ( .ip(n19700), .op(n19739) );
  nand2_1 U16939 ( .ip1(n16410), .ip2(n19739), .op(n15466) );
  nand2_1 U16940 ( .ip1(\pipeline/csr/mbadaddr [8]), .ip2(n16411), .op(n15465)
         );
  nand2_1 U16941 ( .ip1(\pipeline/alu_out_WB [8]), .ip2(n16412), .op(n15464)
         );
  nand2_1 U16942 ( .ip1(n16413), .ip2(\pipeline/PC_WB [8]), .op(n15463) );
  nand4_1 U16943 ( .ip1(n15466), .ip2(n15465), .ip3(n15464), .ip4(n15463), 
        .op(n8692) );
  nand2_1 U16944 ( .ip1(n16368), .ip2(n20400), .op(n15494) );
  nand2_1 U16945 ( .ip1(n16369), .ip2(htif_pcr_req_data[13]), .op(n15493) );
  nand2_1 U16946 ( .ip1(n16335), .ip2(n15467), .op(n15468) );
  nand2_1 U16947 ( .ip1(n16337), .ip2(n15468), .op(n15491) );
  nand2_1 U16948 ( .ip1(ext_interrupts[5]), .ip2(n19599), .op(n15490) );
  nand2_1 U16949 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [13]), .op(
        n15472) );
  nand2_1 U16950 ( .ip1(n16301), .ip2(\pipeline/csr/instret_full [13]), .op(
        n15471) );
  nand2_1 U16951 ( .ip1(n16383), .ip2(\pipeline/csr/from_host [13]), .op(
        n15470) );
  nand2_1 U16952 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [13]), .op(n15469)
         );
  nand4_1 U16953 ( .ip1(n15472), .ip2(n15471), .ip3(n15470), .ip4(n15469), 
        .op(n15476) );
  nand2_1 U16954 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [13]), .op(n15474) );
  nand2_1 U16955 ( .ip1(\pipeline/epc [13]), .ip2(n17305), .op(n15473) );
  nand2_1 U16956 ( .ip1(n15474), .ip2(n15473), .op(n15475) );
  not_ab_or_c_or_d U16957 ( .ip1(n16310), .ip2(\pipeline/csr/mtime_full [45]), 
        .ip3(n15476), .ip4(n15475), .op(n15489) );
  nand2_1 U16958 ( .ip1(\pipeline/csr/mie [13]), .ip2(n18144), .op(n15480) );
  nand2_1 U16959 ( .ip1(n16382), .ip2(\pipeline/csr/mtime_full [13]), .op(
        n15479) );
  nand2_1 U16960 ( .ip1(\pipeline/csr/mtvec [13]), .ip2(n17364), .op(n15478)
         );
  nand2_1 U16961 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [13]), .op(n15477) );
  nand4_1 U16962 ( .ip1(n15480), .ip2(n15479), .ip3(n15478), .ip4(n15477), 
        .op(n15486) );
  nand2_1 U16963 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [45]), .op(
        n15484) );
  nand2_1 U16964 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [13]), .op(
        n15483) );
  nand2_1 U16965 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [45]), .op(
        n15482) );
  nand2_1 U16966 ( .ip1(n16373), .ip2(\pipeline/csr/time_full [45]), .op(
        n15481) );
  nand4_1 U16967 ( .ip1(n15484), .ip2(n15483), .ip3(n15482), .ip4(n15481), 
        .op(n15485) );
  nor2_1 U16968 ( .ip1(n15486), .ip2(n15485), .op(n15488) );
  nand2_1 U16969 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [13]), .op(n15487) );
  nand4_1 U16970 ( .ip1(n15490), .ip2(n15489), .ip3(n15488), .ip4(n15487), 
        .op(n20275) );
  nand2_1 U16971 ( .ip1(n15491), .ip2(n20275), .op(n15492) );
  nand3_1 U16972 ( .ip1(n15494), .ip2(n15493), .ip3(n15492), .op(n22166) );
  nand2_1 U16973 ( .ip1(n16410), .ip2(n22166), .op(n15498) );
  nand2_1 U16974 ( .ip1(\pipeline/csr/mbadaddr [13]), .ip2(n16411), .op(n15497) );
  nand2_1 U16975 ( .ip1(\pipeline/alu_out_WB [13]), .ip2(n16412), .op(n15496)
         );
  nand2_1 U16976 ( .ip1(n16413), .ip2(\pipeline/PC_WB [13]), .op(n15495) );
  nand4_1 U16977 ( .ip1(n15498), .ip2(n15497), .ip3(n15496), .ip4(n15495), 
        .op(n8687) );
  nand2_1 U16978 ( .ip1(n16368), .ip2(n20007), .op(n15526) );
  nand2_1 U16979 ( .ip1(n16369), .ip2(htif_pcr_req_data[17]), .op(n15525) );
  nand2_1 U16980 ( .ip1(n16335), .ip2(n15499), .op(n15500) );
  nand2_1 U16981 ( .ip1(n16337), .ip2(n15500), .op(n15523) );
  nand2_1 U16982 ( .ip1(ext_interrupts[9]), .ip2(n19599), .op(n15522) );
  nand2_1 U16983 ( .ip1(n16373), .ip2(\pipeline/csr/time_full [49]), .op(
        n15504) );
  nand2_1 U16984 ( .ip1(n16301), .ip2(\pipeline/csr/instret_full [17]), .op(
        n15503) );
  nand2_1 U16985 ( .ip1(n16383), .ip2(\pipeline/csr/from_host [17]), .op(
        n15502) );
  nand2_1 U16986 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [17]), .op(n15501)
         );
  nand4_1 U16987 ( .ip1(n15504), .ip2(n15503), .ip3(n15502), .ip4(n15501), 
        .op(n15508) );
  nand2_1 U16988 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [17]), .op(n15506) );
  nand2_1 U16989 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [17]), .op(n15505) );
  nand2_1 U16990 ( .ip1(n15506), .ip2(n15505), .op(n15507) );
  not_ab_or_c_or_d U16991 ( .ip1(n16310), .ip2(\pipeline/csr/mtime_full [49]), 
        .ip3(n15508), .ip4(n15507), .op(n15521) );
  nand2_1 U16992 ( .ip1(\pipeline/csr/mtvec [17]), .ip2(n17364), .op(n15512)
         );
  nand2_1 U16993 ( .ip1(n16382), .ip2(\pipeline/csr/mtime_full [17]), .op(
        n15511) );
  nand2_1 U16994 ( .ip1(\pipeline/csr/mie [17]), .ip2(n18144), .op(n15510) );
  nand2_1 U16995 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [17]), .op(n15509) );
  nand4_1 U16996 ( .ip1(n15512), .ip2(n15511), .ip3(n15510), .ip4(n15509), 
        .op(n15518) );
  nand2_1 U16997 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [49]), .op(
        n15516) );
  nand2_1 U16998 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [17]), .op(
        n15515) );
  nand2_1 U16999 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [49]), .op(
        n15514) );
  nand2_1 U17000 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [17]), .op(
        n15513) );
  nand4_1 U17001 ( .ip1(n15516), .ip2(n15515), .ip3(n15514), .ip4(n15513), 
        .op(n15517) );
  nor2_1 U17002 ( .ip1(n15518), .ip2(n15517), .op(n15520) );
  nand2_1 U17003 ( .ip1(\pipeline/epc [17]), .ip2(n17305), .op(n15519) );
  nand4_1 U17004 ( .ip1(n15522), .ip2(n15521), .ip3(n15520), .ip4(n15519), 
        .op(n20004) );
  nand2_1 U17005 ( .ip1(n15523), .ip2(n20004), .op(n15524) );
  nand3_1 U17006 ( .ip1(n15526), .ip2(n15525), .ip3(n15524), .op(n22183) );
  nand2_1 U17007 ( .ip1(n16410), .ip2(n22183), .op(n15530) );
  nand2_1 U17008 ( .ip1(\pipeline/csr/mbadaddr [17]), .ip2(n16411), .op(n15529) );
  nand2_1 U17009 ( .ip1(\pipeline/alu_out_WB [17]), .ip2(n16412), .op(n15528)
         );
  nand2_1 U17010 ( .ip1(n16413), .ip2(\pipeline/PC_WB [17]), .op(n15527) );
  nand4_1 U17011 ( .ip1(n15530), .ip2(n15529), .ip3(n15528), .ip4(n15527), 
        .op(n8683) );
  nand2_1 U17012 ( .ip1(n16368), .ip2(n20586), .op(n15560) );
  nand2_1 U17013 ( .ip1(n16369), .ip2(htif_pcr_req_data[21]), .op(n15559) );
  nand2_1 U17014 ( .ip1(n16335), .ip2(n15531), .op(n15532) );
  nand2_1 U17015 ( .ip1(n16337), .ip2(n15532), .op(n15557) );
  inv_1 U17016 ( .ip(\pipeline/epc [21]), .op(n18638) );
  inv_1 U17017 ( .ip(n17305), .op(n15869) );
  nor2_1 U17018 ( .ip1(n18638), .ip2(n15869), .op(n15546) );
  inv_1 U17019 ( .ip(\pipeline/csr/mtimecmp [21]), .op(n22370) );
  nor2_1 U17020 ( .ip1(n22370), .ip2(n15533), .op(n15537) );
  nand2_1 U17021 ( .ip1(\pipeline/csr/mie [21]), .ip2(n18144), .op(n15535) );
  nand2_1 U17022 ( .ip1(n16382), .ip2(\pipeline/csr/mtime_full [21]), .op(
        n15534) );
  nand2_1 U17023 ( .ip1(n15535), .ip2(n15534), .op(n15536) );
  not_ab_or_c_or_d U17024 ( .ip1(n17364), .ip2(\pipeline/csr/mtvec [21]), 
        .ip3(n15537), .ip4(n15536), .op(n15544) );
  inv_1 U17025 ( .ip(\pipeline/csr/time_full [21]), .op(n17643) );
  nor2_1 U17026 ( .ip1(n15538), .ip2(n17643), .op(n15540) );
  inv_1 U17027 ( .ip(n16373), .op(n15864) );
  inv_1 U17028 ( .ip(\pipeline/csr/time_full [53]), .op(n17649) );
  nor2_1 U17029 ( .ip1(n15864), .ip2(n17649), .op(n15539) );
  nor2_1 U17030 ( .ip1(n15540), .ip2(n15539), .op(n15543) );
  nand2_1 U17031 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [21]), .op(
        n15542) );
  nand2_1 U17032 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [53]), .op(
        n15541) );
  nand4_1 U17033 ( .ip1(n15544), .ip2(n15543), .ip3(n15542), .ip4(n15541), 
        .op(n15545) );
  not_ab_or_c_or_d U17034 ( .ip1(n19599), .ip2(ext_interrupts[13]), .ip3(
        n15546), .ip4(n15545), .op(n15556) );
  nand2_1 U17035 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [53]), .op(
        n15550) );
  nand2_1 U17036 ( .ip1(n16301), .ip2(\pipeline/csr/instret_full [21]), .op(
        n15549) );
  nand2_1 U17037 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [21]), .op(n15548)
         );
  nand2_1 U17038 ( .ip1(n16383), .ip2(\pipeline/csr/from_host [21]), .op(
        n15547) );
  nand4_1 U17039 ( .ip1(n15550), .ip2(n15549), .ip3(n15548), .ip4(n15547), 
        .op(n15554) );
  nand2_1 U17040 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [21]), .op(n15552) );
  nand2_1 U17041 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [21]), .op(n15551) );
  nand2_1 U17042 ( .ip1(n15552), .ip2(n15551), .op(n15553) );
  not_ab_or_c_or_d U17043 ( .ip1(n16310), .ip2(\pipeline/csr/mtime_full [53]), 
        .ip3(n15554), .ip4(n15553), .op(n15555) );
  nand2_1 U17044 ( .ip1(n15556), .ip2(n15555), .op(n20469) );
  nand2_1 U17045 ( .ip1(n15557), .ip2(n20469), .op(n15558) );
  nand3_1 U17046 ( .ip1(n15560), .ip2(n15559), .ip3(n15558), .op(n22368) );
  nand2_1 U17047 ( .ip1(n16410), .ip2(n22368), .op(n15564) );
  nand2_1 U17048 ( .ip1(\pipeline/csr/mbadaddr [21]), .ip2(n16411), .op(n15563) );
  nand2_1 U17049 ( .ip1(\pipeline/alu_out_WB [21]), .ip2(n16412), .op(n15562)
         );
  nand2_1 U17050 ( .ip1(n16413), .ip2(\pipeline/PC_WB [21]), .op(n15561) );
  nand4_1 U17051 ( .ip1(n15564), .ip2(n15563), .ip3(n15562), .ip4(n15561), 
        .op(n8679) );
  nand2_1 U17052 ( .ip1(n16368), .ip2(n15565), .op(n15592) );
  nand2_1 U17053 ( .ip1(n16369), .ip2(htif_pcr_req_data[25]), .op(n15591) );
  nand2_1 U17054 ( .ip1(n16335), .ip2(n20158), .op(n15566) );
  nand2_1 U17055 ( .ip1(n16337), .ip2(n15566), .op(n15589) );
  nand2_1 U17056 ( .ip1(ext_interrupts[17]), .ip2(n19599), .op(n15588) );
  nand2_1 U17057 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [25]), .op(
        n15570) );
  nand2_1 U17058 ( .ip1(n16301), .ip2(\pipeline/csr/instret_full [25]), .op(
        n15569) );
  nand2_1 U17059 ( .ip1(n16383), .ip2(\pipeline/csr/from_host [25]), .op(
        n15568) );
  nand2_1 U17060 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [25]), .op(n15567)
         );
  nand4_1 U17061 ( .ip1(n15570), .ip2(n15569), .ip3(n15568), .ip4(n15567), 
        .op(n15574) );
  nand2_1 U17062 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [25]), .op(n15572) );
  nand2_1 U17063 ( .ip1(\pipeline/epc [25]), .ip2(n17305), .op(n15571) );
  nand2_1 U17064 ( .ip1(n15572), .ip2(n15571), .op(n15573) );
  not_ab_or_c_or_d U17065 ( .ip1(n16310), .ip2(\pipeline/csr/mtime_full [57]), 
        .ip3(n15574), .ip4(n15573), .op(n15587) );
  nand2_1 U17066 ( .ip1(n16382), .ip2(\pipeline/csr/mtime_full [25]), .op(
        n15578) );
  nand2_1 U17067 ( .ip1(\pipeline/csr/mtvec [25]), .ip2(n17364), .op(n15577)
         );
  nand2_1 U17068 ( .ip1(\pipeline/csr/mie [25]), .ip2(n18144), .op(n15576) );
  nand2_1 U17069 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [25]), .op(n15575) );
  nand4_1 U17070 ( .ip1(n15578), .ip2(n15577), .ip3(n15576), .ip4(n15575), 
        .op(n15584) );
  nand2_1 U17071 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [57]), .op(
        n15582) );
  nand2_1 U17072 ( .ip1(n16373), .ip2(\pipeline/csr/time_full [57]), .op(
        n15581) );
  nand2_1 U17073 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [25]), .op(
        n15580) );
  nand2_1 U17074 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [57]), .op(
        n15579) );
  nand4_1 U17075 ( .ip1(n15582), .ip2(n15581), .ip3(n15580), .ip4(n15579), 
        .op(n15583) );
  nor2_1 U17076 ( .ip1(n15584), .ip2(n15583), .op(n15586) );
  nand2_1 U17077 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [25]), .op(n15585) );
  nand4_1 U17078 ( .ip1(n15588), .ip2(n15587), .ip3(n15586), .ip4(n15585), 
        .op(n20162) );
  nand2_1 U17079 ( .ip1(n15589), .ip2(n20162), .op(n15590) );
  nand3_1 U17080 ( .ip1(n15592), .ip2(n15591), .ip3(n15590), .op(n22217) );
  nand2_1 U17081 ( .ip1(n16410), .ip2(n22217), .op(n15596) );
  nand2_1 U17082 ( .ip1(\pipeline/csr/mbadaddr [25]), .ip2(n16411), .op(n15595) );
  nand2_1 U17083 ( .ip1(\pipeline/alu_out_WB [25]), .ip2(n16412), .op(n15594)
         );
  nand2_1 U17084 ( .ip1(n16413), .ip2(\pipeline/PC_WB [25]), .op(n15593) );
  nand4_1 U17085 ( .ip1(n15596), .ip2(n15595), .ip3(n15594), .ip4(n15593), 
        .op(n8675) );
  nand2_1 U17086 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [50]), .op(
        n15601) );
  nand2_1 U17087 ( .ip1(n16301), .ip2(\pipeline/csr/instret_full [18]), .op(
        n15600) );
  nand2_1 U17088 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [18]), .op(n15599)
         );
  nand2_1 U17089 ( .ip1(n16383), .ip2(\pipeline/csr/from_host [18]), .op(
        n15598) );
  nand4_1 U17090 ( .ip1(n15601), .ip2(n15600), .ip3(n15599), .ip4(n15598), 
        .op(n15605) );
  nand2_1 U17091 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [18]), .op(n15603) );
  nand2_1 U17092 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [18]), .op(n15602) );
  nand2_1 U17093 ( .ip1(n15603), .ip2(n15602), .op(n15604) );
  not_ab_or_c_or_d U17094 ( .ip1(n16310), .ip2(\pipeline/csr/mtime_full [50]), 
        .ip3(n15605), .ip4(n15604), .op(n15619) );
  nand2_1 U17095 ( .ip1(\pipeline/csr/mie [18]), .ip2(n18144), .op(n15609) );
  nand2_1 U17096 ( .ip1(n16382), .ip2(\pipeline/csr/mtime_full [18]), .op(
        n15608) );
  nand2_1 U17097 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [18]), .op(n15607) );
  nand2_1 U17098 ( .ip1(\pipeline/csr/mtvec [18]), .ip2(n17364), .op(n15606)
         );
  nand4_1 U17099 ( .ip1(n15609), .ip2(n15608), .ip3(n15607), .ip4(n15606), 
        .op(n15615) );
  nand2_1 U17100 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [50]), .op(
        n15613) );
  nand2_1 U17101 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [18]), .op(
        n15612) );
  nand2_1 U17102 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [18]), .op(
        n15611) );
  nand2_1 U17103 ( .ip1(n16373), .ip2(\pipeline/csr/time_full [50]), .op(
        n15610) );
  nand4_1 U17104 ( .ip1(n15613), .ip2(n15612), .ip3(n15611), .ip4(n15610), 
        .op(n15614) );
  nor2_1 U17105 ( .ip1(n15615), .ip2(n15614), .op(n15618) );
  nand2_1 U17106 ( .ip1(\pipeline/epc [18]), .ip2(n17305), .op(n15617) );
  nand2_1 U17107 ( .ip1(ext_interrupts[10]), .ip2(n19599), .op(n15616) );
  and4_1 U17108 ( .ip1(n15619), .ip2(n15618), .ip3(n15617), .ip4(n15616), .op(
        n20017) );
  nor2_1 U17109 ( .ip1(n15597), .ip2(n16401), .op(n15620) );
  nor2_1 U17110 ( .ip1(n15620), .ip2(n16403), .op(n15621) );
  nor2_1 U17111 ( .ip1(n20017), .ip2(n15621), .op(n15623) );
  and2_1 U17112 ( .ip1(n16369), .ip2(htif_pcr_req_data[18]), .op(n15622) );
  not_ab_or_c_or_d U17113 ( .ip1(n16368), .ip2(n15597), .ip3(n15623), .ip4(
        n15622), .op(n18572) );
  inv_1 U17114 ( .ip(n18572), .op(n18563) );
  nand2_1 U17115 ( .ip1(n16410), .ip2(n18563), .op(n15627) );
  nand2_1 U17116 ( .ip1(n16413), .ip2(\pipeline/PC_WB [18]), .op(n15626) );
  nand2_1 U17117 ( .ip1(\pipeline/csr/mbadaddr [18]), .ip2(n16411), .op(n15625) );
  nand2_1 U17118 ( .ip1(\pipeline/alu_out_WB [18]), .ip2(n16412), .op(n15624)
         );
  nand4_1 U17119 ( .ip1(n15627), .ip2(n15626), .ip3(n15625), .ip4(n15624), 
        .op(n8682) );
  nand2_1 U17120 ( .ip1(n15628), .ip2(n16368), .op(n15655) );
  nand2_1 U17121 ( .ip1(n16369), .ip2(htif_pcr_req_data[19]), .op(n15654) );
  nand2_1 U17122 ( .ip1(n16335), .ip2(n20571), .op(n15629) );
  nand2_1 U17123 ( .ip1(n16337), .ip2(n15629), .op(n15652) );
  nand2_1 U17124 ( .ip1(ext_interrupts[11]), .ip2(n19599), .op(n15651) );
  nand2_1 U17125 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [51]), .op(
        n15633) );
  nand2_1 U17126 ( .ip1(n16301), .ip2(\pipeline/csr/instret_full [19]), .op(
        n15632) );
  nand2_1 U17127 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [19]), .op(n15631)
         );
  nand2_1 U17128 ( .ip1(n16383), .ip2(\pipeline/csr/from_host [19]), .op(
        n15630) );
  nand4_1 U17129 ( .ip1(n15633), .ip2(n15632), .ip3(n15631), .ip4(n15630), 
        .op(n15637) );
  nand2_1 U17130 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [19]), .op(n15635) );
  nand2_1 U17131 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [19]), .op(n15634) );
  nand2_1 U17132 ( .ip1(n15635), .ip2(n15634), .op(n15636) );
  not_ab_or_c_or_d U17133 ( .ip1(n16310), .ip2(\pipeline/csr/mtime_full [51]), 
        .ip3(n15637), .ip4(n15636), .op(n15650) );
  nand2_1 U17134 ( .ip1(\pipeline/csr/mie [19]), .ip2(n18144), .op(n15641) );
  nand2_1 U17135 ( .ip1(n16382), .ip2(\pipeline/csr/mtime_full [19]), .op(
        n15640) );
  nand2_1 U17136 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [19]), .op(n15639) );
  nand2_1 U17137 ( .ip1(\pipeline/csr/mtvec [19]), .ip2(n17364), .op(n15638)
         );
  nand4_1 U17138 ( .ip1(n15641), .ip2(n15640), .ip3(n15639), .ip4(n15638), 
        .op(n15647) );
  nand2_1 U17139 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [51]), .op(
        n15645) );
  nand2_1 U17140 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [19]), .op(
        n15644) );
  nand2_1 U17141 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [19]), .op(
        n15643) );
  nand2_1 U17142 ( .ip1(n16373), .ip2(\pipeline/csr/time_full [51]), .op(
        n15642) );
  nand4_1 U17143 ( .ip1(n15645), .ip2(n15644), .ip3(n15643), .ip4(n15642), 
        .op(n15646) );
  nor2_1 U17144 ( .ip1(n15647), .ip2(n15646), .op(n15649) );
  nand2_1 U17145 ( .ip1(\pipeline/epc [19]), .ip2(n17305), .op(n15648) );
  nand4_1 U17146 ( .ip1(n15651), .ip2(n15650), .ip3(n15649), .ip4(n15648), 
        .op(n20563) );
  nand2_1 U17147 ( .ip1(n15652), .ip2(n20563), .op(n15653) );
  nand3_1 U17148 ( .ip1(n15655), .ip2(n15654), .ip3(n15653), .op(n22189) );
  nand2_1 U17149 ( .ip1(n16410), .ip2(n22189), .op(n15659) );
  nand2_1 U17150 ( .ip1(\pipeline/csr/mbadaddr [19]), .ip2(n16411), .op(n15658) );
  nand2_1 U17151 ( .ip1(\pipeline/alu_out_WB [19]), .ip2(n16412), .op(n15657)
         );
  nand2_1 U17152 ( .ip1(n16413), .ip2(\pipeline/PC_WB [19]), .op(n15656) );
  nand4_1 U17153 ( .ip1(n15659), .ip2(n15658), .ip3(n15657), .ip4(n15656), 
        .op(n8681) );
  mux2_1 U17154 ( .ip1(n15661), .ip2(n15660), .s(\pipeline/dmem_type[2] ), 
        .op(n15687) );
  nand2_1 U17155 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [4]), .op(
        n15665) );
  nand2_1 U17156 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [4]), .op(n15664) );
  nand2_1 U17157 ( .ip1(n16373), .ip2(\pipeline/csr/time_full [36]), .op(
        n15663) );
  nand2_1 U17158 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [36]), .op(
        n15662) );
  and4_1 U17159 ( .ip1(n15665), .ip2(n15664), .ip3(n15663), .ip4(n15662), .op(
        n15684) );
  inv_1 U17160 ( .ip(\pipeline/epc [4]), .op(n17966) );
  nor2_1 U17161 ( .ip1(n17966), .ip2(n15869), .op(n15680) );
  inv_1 U17162 ( .ip(\pipeline/csr/instret_full [4]), .op(n21009) );
  nor2_1 U17163 ( .ip1(n16380), .ip2(n21009), .op(n15668) );
  inv_1 U17164 ( .ip(n16383), .op(n17833) );
  inv_1 U17165 ( .ip(\pipeline/csr/from_host [4]), .op(n15666) );
  nor2_1 U17166 ( .ip1(n17833), .ip2(n15666), .op(n15667) );
  not_ab_or_c_or_d U17167 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [4]), 
        .ip3(n15668), .ip4(n15667), .op(n15678) );
  nand2_1 U17168 ( .ip1(n18144), .ip2(\pipeline/csr/mie [4]), .op(n15672) );
  nand2_1 U17169 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [4]), .op(n15671)
         );
  nand2_1 U17170 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [36]), .op(
        n15670) );
  nand2_1 U17171 ( .ip1(\pipeline/csr/mtvec [4]), .ip2(n17364), .op(n15669) );
  and4_1 U17172 ( .ip1(n15672), .ip2(n15671), .ip3(n15670), .ip4(n15669), .op(
        n15677) );
  nand2_1 U17173 ( .ip1(n16382), .ip2(\pipeline/csr/mtime_full [4]), .op(
        n15676) );
  nor2_1 U17174 ( .ip1(n15674), .ip2(n15673), .op(n20964) );
  nand2_1 U17175 ( .ip1(n20964), .ip2(\pipeline/csr/priv_stack [4]), .op(
        n15675) );
  nand4_1 U17176 ( .ip1(n15678), .ip2(n15677), .ip3(n15676), .ip4(n15675), 
        .op(n15679) );
  not_ab_or_c_or_d U17177 ( .ip1(\pipeline/csr/mbadaddr [4]), .ip2(n16396), 
        .ip3(n15680), .ip4(n15679), .op(n15683) );
  nand2_1 U17178 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [4]), .op(n15682)
         );
  nand2_1 U17179 ( .ip1(n16310), .ip2(\pipeline/csr/mtime_full [36]), .op(
        n15681) );
  nand4_1 U17180 ( .ip1(n15684), .ip2(n15683), .ip3(n15682), .ip4(n15681), 
        .op(n21028) );
  nand3_1 U17181 ( .ip1(n15687), .ip2(n16335), .ip3(n21028), .op(n15686) );
  nand2_1 U17182 ( .ip1(n16369), .ip2(htif_pcr_req_data[4]), .op(n15685) );
  and2_1 U17183 ( .ip1(n15686), .ip2(n15685), .op(n17951) );
  inv_1 U17184 ( .ip(n16019), .op(n16073) );
  inv_1 U17185 ( .ip(n15687), .op(n17948) );
  nand2_1 U17186 ( .ip1(n16073), .ip2(n17948), .op(n15688) );
  nand2_1 U17187 ( .ip1(n17951), .ip2(n15688), .op(n17972) );
  nand2_1 U17188 ( .ip1(n16410), .ip2(n17972), .op(n15692) );
  nand2_1 U17189 ( .ip1(n16413), .ip2(\pipeline/PC_WB [4]), .op(n15691) );
  nand2_1 U17190 ( .ip1(n16411), .ip2(\pipeline/csr/mbadaddr [4]), .op(n15690)
         );
  nand2_1 U17191 ( .ip1(\pipeline/alu_out_WB [4]), .ip2(n16412), .op(n15689)
         );
  nand4_1 U17192 ( .ip1(n15692), .ip2(n15691), .ip3(n15690), .ip4(n15689), 
        .op(n8696) );
  nand2_1 U17193 ( .ip1(n16368), .ip2(n15693), .op(n15720) );
  nand2_1 U17194 ( .ip1(n16369), .ip2(htif_pcr_req_data[14]), .op(n15719) );
  nand2_1 U17195 ( .ip1(n16335), .ip2(n20424), .op(n15694) );
  nand2_1 U17196 ( .ip1(n16337), .ip2(n15694), .op(n15717) );
  nand2_1 U17197 ( .ip1(ext_interrupts[6]), .ip2(n19599), .op(n15716) );
  nand2_1 U17198 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [46]), .op(
        n15698) );
  nand2_1 U17199 ( .ip1(n16301), .ip2(\pipeline/csr/instret_full [14]), .op(
        n15697) );
  nand2_1 U17200 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [14]), .op(n15696)
         );
  nand2_1 U17201 ( .ip1(n16383), .ip2(\pipeline/csr/from_host [14]), .op(
        n15695) );
  nand4_1 U17202 ( .ip1(n15698), .ip2(n15697), .ip3(n15696), .ip4(n15695), 
        .op(n15702) );
  nand2_1 U17203 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [14]), .op(n15700) );
  nand2_1 U17204 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [14]), .op(n15699) );
  nand2_1 U17205 ( .ip1(n15700), .ip2(n15699), .op(n15701) );
  not_ab_or_c_or_d U17206 ( .ip1(n16310), .ip2(\pipeline/csr/mtime_full [46]), 
        .ip3(n15702), .ip4(n15701), .op(n15715) );
  nand2_1 U17207 ( .ip1(\pipeline/csr/mie [14]), .ip2(n18144), .op(n15706) );
  nand2_1 U17208 ( .ip1(n16382), .ip2(\pipeline/csr/mtime_full [14]), .op(
        n15705) );
  nand2_1 U17209 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [14]), .op(n15704) );
  nand2_1 U17210 ( .ip1(\pipeline/csr/mtvec [14]), .ip2(n17364), .op(n15703)
         );
  nand4_1 U17211 ( .ip1(n15706), .ip2(n15705), .ip3(n15704), .ip4(n15703), 
        .op(n15712) );
  nand2_1 U17212 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [46]), .op(
        n15710) );
  nand2_1 U17213 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [14]), .op(
        n15709) );
  nand2_1 U17214 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [14]), .op(
        n15708) );
  nand2_1 U17215 ( .ip1(n16373), .ip2(\pipeline/csr/time_full [46]), .op(
        n15707) );
  nand4_1 U17216 ( .ip1(n15710), .ip2(n15709), .ip3(n15708), .ip4(n15707), 
        .op(n15711) );
  nor2_1 U17217 ( .ip1(n15712), .ip2(n15711), .op(n15714) );
  nand2_1 U17218 ( .ip1(\pipeline/epc [14]), .ip2(n17305), .op(n15713) );
  nand4_1 U17219 ( .ip1(n15716), .ip2(n15715), .ip3(n15714), .ip4(n15713), 
        .op(n19892) );
  nand2_1 U17220 ( .ip1(n15717), .ip2(n19892), .op(n15718) );
  nand3_1 U17221 ( .ip1(n15720), .ip2(n15719), .ip3(n15718), .op(n22171) );
  nand2_1 U17222 ( .ip1(n16410), .ip2(n22171), .op(n15724) );
  nand2_1 U17223 ( .ip1(\pipeline/csr/mbadaddr [14]), .ip2(n16411), .op(n15723) );
  nand2_1 U17224 ( .ip1(\pipeline/alu_out_WB [14]), .ip2(n16412), .op(n15722)
         );
  nand2_1 U17225 ( .ip1(n16413), .ip2(\pipeline/PC_WB [14]), .op(n15721) );
  nand4_1 U17226 ( .ip1(n15724), .ip2(n15723), .ip3(n15722), .ip4(n15721), 
        .op(n8686) );
  nand2_1 U17227 ( .ip1(n16480), .ip2(n22896), .op(n15960) );
  nor2_1 U17228 ( .ip1(n15726), .ip2(n15960), .op(n15753) );
  nand2_1 U17229 ( .ip1(n17765), .ip2(n15725), .op(n15961) );
  nor2_1 U17230 ( .ip1(n15726), .ip2(n15961), .op(n15751) );
  nand2_1 U17231 ( .ip1(n16310), .ip2(\pipeline/csr/mtime_full [47]), .op(
        n15730) );
  nand2_1 U17232 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [15]), .op(n15729) );
  nand2_1 U17233 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [15]), .op(n15728) );
  nand2_1 U17234 ( .ip1(\pipeline/epc [15]), .ip2(n17305), .op(n15727) );
  nand4_1 U17235 ( .ip1(n15730), .ip2(n15729), .ip3(n15728), .ip4(n15727), 
        .op(n15749) );
  inv_1 U17236 ( .ip(\pipeline/csr/mtime_full [15]), .op(n19611) );
  nor2_1 U17237 ( .ip1(n15971), .ip2(n19611), .op(n15733) );
  nor2_1 U17238 ( .ip1(n15731), .ip2(n22100), .op(n15732) );
  not_ab_or_c_or_d U17239 ( .ip1(n16383), .ip2(\pipeline/csr/from_host [15]), 
        .ip3(n15733), .ip4(n15732), .op(n15737) );
  nand2_1 U17240 ( .ip1(ext_interrupts[7]), .ip2(n19599), .op(n15736) );
  nand2_1 U17241 ( .ip1(n16301), .ip2(\pipeline/csr/instret_full [15]), .op(
        n15735) );
  nand2_1 U17242 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [15]), .op(n15734)
         );
  nand4_1 U17243 ( .ip1(n15737), .ip2(n15736), .ip3(n15735), .ip4(n15734), 
        .op(n15748) );
  nand2_1 U17244 ( .ip1(\pipeline/csr/mie [15]), .ip2(n18144), .op(n15741) );
  nand2_1 U17245 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [15]), .op(n15740) );
  nand2_1 U17246 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [47]), .op(
        n15739) );
  nand2_1 U17247 ( .ip1(\pipeline/csr/mtvec [15]), .ip2(n17364), .op(n15738)
         );
  nand4_1 U17248 ( .ip1(n15741), .ip2(n15740), .ip3(n15739), .ip4(n15738), 
        .op(n15747) );
  nand2_1 U17249 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [15]), .op(
        n15745) );
  nand2_1 U17250 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [47]), .op(
        n15744) );
  nand2_1 U17251 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [15]), .op(
        n15743) );
  nand2_1 U17252 ( .ip1(n16373), .ip2(\pipeline/csr/time_full [47]), .op(
        n15742) );
  nand4_1 U17253 ( .ip1(n15745), .ip2(n15744), .ip3(n15743), .ip4(n15742), 
        .op(n15746) );
  nor4_1 U17254 ( .ip1(n15749), .ip2(n15748), .ip3(n15747), .ip4(n15746), .op(
        n19487) );
  nor2_1 U17255 ( .ip1(n19487), .ip2(n16401), .op(n15750) );
  nor2_1 U17256 ( .ip1(n15751), .ip2(n15750), .op(n15752) );
  or2_1 U17257 ( .ip1(n15753), .ip2(n15752), .op(n15755) );
  nand2_1 U17258 ( .ip1(n16369), .ip2(htif_pcr_req_data[15]), .op(n15754) );
  nand2_1 U17259 ( .ip1(n15755), .ip2(n15754), .op(n22177) );
  nand2_1 U17260 ( .ip1(n16410), .ip2(n22177), .op(n15759) );
  nand2_1 U17261 ( .ip1(n16411), .ip2(\pipeline/csr/mbadaddr [15]), .op(n15758) );
  nand2_1 U17262 ( .ip1(\pipeline/alu_out_WB [15]), .ip2(n16412), .op(n15757)
         );
  nand2_1 U17263 ( .ip1(n16413), .ip2(\pipeline/PC_WB [15]), .op(n15756) );
  nand4_1 U17264 ( .ip1(n15759), .ip2(n15758), .ip3(n15757), .ip4(n15756), 
        .op(n8685) );
  nand2_1 U17265 ( .ip1(n16310), .ip2(\pipeline/csr/mtime_full [34]), .op(
        n15763) );
  nand2_1 U17266 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [2]), .op(n15762)
         );
  nor2_1 U17267 ( .ip1(n22093), .ip2(n22110), .op(n16039) );
  nand2_1 U17268 ( .ip1(n16039), .ip2(\pipeline/csr/mecode [2]), .op(n15761)
         );
  nand2_1 U17269 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [2]), .op(n15760)
         );
  nand4_1 U17270 ( .ip1(n15763), .ip2(n15762), .ip3(n15761), .ip4(n15760), 
        .op(n15781) );
  and2_1 U17271 ( .ip1(n16383), .ip2(\pipeline/csr/from_host [2]), .op(n15765)
         );
  inv_1 U17272 ( .ip(\pipeline/csr/instret_full [2]), .op(n20998) );
  nor2_1 U17273 ( .ip1(n16380), .ip2(n20998), .op(n15764) );
  not_ab_or_c_or_d U17274 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [2]), 
        .ip3(n15765), .ip4(n15764), .op(n15769) );
  nand2_1 U17275 ( .ip1(\pipeline/epc [2]), .ip2(n17305), .op(n15768) );
  nand2_1 U17276 ( .ip1(\pipeline/prv [1]), .ip2(n20964), .op(n15767) );
  nand2_1 U17277 ( .ip1(n16382), .ip2(\pipeline/csr/mtime_full [2]), .op(
        n15766) );
  nand4_1 U17278 ( .ip1(n15769), .ip2(n15768), .ip3(n15767), .ip4(n15766), 
        .op(n15780) );
  nand2_1 U17279 ( .ip1(n18144), .ip2(\pipeline/csr/mie [2]), .op(n15773) );
  nand2_1 U17280 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [2]), .op(n15772)
         );
  nand2_1 U17281 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [34]), .op(
        n15771) );
  nand2_1 U17282 ( .ip1(\pipeline/csr/mtvec [2]), .ip2(n17364), .op(n15770) );
  nand4_1 U17283 ( .ip1(n15773), .ip2(n15772), .ip3(n15771), .ip4(n15770), 
        .op(n15779) );
  nand2_1 U17284 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [2]), .op(
        n15777) );
  nand2_1 U17285 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [2]), .op(n15776) );
  nand2_1 U17286 ( .ip1(n16373), .ip2(\pipeline/csr/time_full [34]), .op(
        n15775) );
  nand2_1 U17287 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [34]), .op(
        n15774) );
  nand4_1 U17288 ( .ip1(n15777), .ip2(n15776), .ip3(n15775), .ip4(n15774), 
        .op(n15778) );
  or4_1 U17289 ( .ip1(n15781), .ip2(n15780), .ip3(n15779), .ip4(n15778), .op(
        n21150) );
  nand2_1 U17290 ( .ip1(n16403), .ip2(n15782), .op(n15785) );
  nor2_1 U17291 ( .ip1(\pipeline/dmem_type[2] ), .ip2(n15789), .op(n15783) );
  nand2_1 U17292 ( .ip1(n16335), .ip2(n15783), .op(n15784) );
  nand2_1 U17293 ( .ip1(n15785), .ip2(n15784), .op(n15788) );
  and2_1 U17294 ( .ip1(n16369), .ip2(htif_pcr_req_data[2]), .op(n15787) );
  and3_1 U17295 ( .ip1(n17949), .ip2(\pipeline/inst_DX [17]), .ip3(
        \pipeline/dmem_type[2] ), .op(n15786) );
  not_ab_or_c_or_d U17296 ( .ip1(n21150), .ip2(n15788), .ip3(n15787), .ip4(
        n15786), .op(n15791) );
  nand2_1 U17297 ( .ip1(n16368), .ip2(n15789), .op(n15790) );
  nand2_1 U17298 ( .ip1(n15791), .ip2(n15790), .op(n22351) );
  nand2_1 U17299 ( .ip1(n16410), .ip2(n22351), .op(n15795) );
  nand2_1 U17300 ( .ip1(\pipeline/csr/mbadaddr [2]), .ip2(n16411), .op(n15794)
         );
  nand2_1 U17301 ( .ip1(\pipeline/alu_out_WB [2]), .ip2(n16412), .op(n15793)
         );
  nand2_1 U17302 ( .ip1(n16413), .ip2(\pipeline/PC_WB [2]), .op(n15792) );
  nand4_1 U17303 ( .ip1(n15795), .ip2(n15794), .ip3(n15793), .ip4(n15792), 
        .op(n8698) );
  nand2_1 U17304 ( .ip1(n16368), .ip2(n15796), .op(n15828) );
  nand2_1 U17305 ( .ip1(n16039), .ip2(\pipeline/csr/mecode [3]), .op(n15800)
         );
  nand2_1 U17306 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [3]), .op(n15799)
         );
  nand2_1 U17307 ( .ip1(\pipeline/csr/mip_3 ), .ip2(n19599), .op(n15798) );
  nand2_1 U17308 ( .ip1(\pipeline/epc [3]), .ip2(n17305), .op(n15797) );
  and4_1 U17309 ( .ip1(n15800), .ip2(n15799), .ip3(n15798), .ip4(n15797), .op(
        n15820) );
  inv_1 U17310 ( .ip(\pipeline/csr/mtime_full [3]), .op(n21191) );
  nor2_1 U17311 ( .ip1(n15971), .ip2(n21191), .op(n15805) );
  nand2_1 U17312 ( .ip1(n16301), .ip2(\pipeline/csr/instret_full [3]), .op(
        n15803) );
  nand2_1 U17313 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [3]), .op(n15802)
         );
  nand2_1 U17314 ( .ip1(n16383), .ip2(\pipeline/csr/from_host [3]), .op(n15801) );
  nand3_1 U17315 ( .ip1(n15803), .ip2(n15802), .ip3(n15801), .op(n15804) );
  not_ab_or_c_or_d U17316 ( .ip1(n20964), .ip2(\pipeline/csr/priv_stack [3]), 
        .ip3(n15805), .ip4(n15804), .op(n15819) );
  nand2_1 U17317 ( .ip1(\pipeline/csr/mie [3]), .ip2(n18144), .op(n15809) );
  nand2_1 U17318 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [3]), .op(n15808)
         );
  nand2_1 U17319 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [35]), .op(
        n15807) );
  nand2_1 U17320 ( .ip1(\pipeline/csr/mtvec [3]), .ip2(n17364), .op(n15806) );
  and4_1 U17321 ( .ip1(n15809), .ip2(n15808), .ip3(n15807), .ip4(n15806), .op(
        n15818) );
  inv_1 U17322 ( .ip(\pipeline/csr/mtime_full [35]), .op(n15810) );
  nor2_1 U17323 ( .ip1(n16338), .ip2(n15810), .op(n15816) );
  nand2_1 U17324 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [3]), .op(
        n15814) );
  nand2_1 U17325 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [3]), .op(n15813) );
  nand2_1 U17326 ( .ip1(n16373), .ip2(\pipeline/csr/time_full [35]), .op(
        n15812) );
  nand2_1 U17327 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [35]), .op(
        n15811) );
  nand4_1 U17328 ( .ip1(n15814), .ip2(n15813), .ip3(n15812), .ip4(n15811), 
        .op(n15815) );
  not_ab_or_c_or_d U17329 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [3]), 
        .ip3(n15816), .ip4(n15815), .op(n15817) );
  nand4_1 U17330 ( .ip1(n15820), .ip2(n15819), .ip3(n15818), .ip4(n15817), 
        .op(n17882) );
  nand3_1 U17331 ( .ip1(n17855), .ip2(n16335), .ip3(n17765), .op(n15823) );
  nand2_1 U17332 ( .ip1(n16403), .ip2(n15821), .op(n15822) );
  nand2_1 U17333 ( .ip1(n15823), .ip2(n15822), .op(n15824) );
  nand2_1 U17334 ( .ip1(n17882), .ip2(n15824), .op(n15827) );
  nand2_1 U17335 ( .ip1(n16369), .ip2(htif_pcr_req_data[3]), .op(n15826) );
  nand3_1 U17336 ( .ip1(\pipeline/inst_DX [18]), .ip2(\pipeline/dmem_type[2] ), 
        .ip3(n17949), .op(n15825) );
  nand4_1 U17337 ( .ip1(n15828), .ip2(n15827), .ip3(n15826), .ip4(n15825), 
        .op(n21223) );
  nand2_1 U17338 ( .ip1(n16410), .ip2(n21223), .op(n15832) );
  nand2_1 U17339 ( .ip1(\pipeline/csr/mbadaddr [3]), .ip2(n16411), .op(n15831)
         );
  nand2_1 U17340 ( .ip1(\pipeline/alu_out_WB [3]), .ip2(n16412), .op(n15830)
         );
  nand2_1 U17341 ( .ip1(n16413), .ip2(\pipeline/PC_WB [3]), .op(n15829) );
  nand4_1 U17342 ( .ip1(n15832), .ip2(n15831), .ip3(n15830), .ip4(n15829), 
        .op(n8697) );
  mux2_1 U17343 ( .ip1(n17334), .ip2(n15833), .s(\pipeline/dmem_type[2] ), 
        .op(n16062) );
  nor2_1 U17344 ( .ip1(n16062), .ip2(n16019), .op(n15856) );
  nand2_1 U17345 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [33]), .op(
        n15837) );
  nand2_1 U17346 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [1]), .op(
        n15836) );
  nand2_1 U17347 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [33]), .op(
        n15835) );
  nand2_1 U17348 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [1]), .op(n15834) );
  nand4_1 U17349 ( .ip1(n15837), .ip2(n15836), .ip3(n15835), .ip4(n15834), 
        .op(n15843) );
  nand2_1 U17350 ( .ip1(n16373), .ip2(\pipeline/csr/time_full [33]), .op(
        n15841) );
  nand2_1 U17351 ( .ip1(n16301), .ip2(\pipeline/csr/instret_full [1]), .op(
        n15840) );
  nand2_1 U17352 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [1]), .op(n15839)
         );
  nand2_1 U17353 ( .ip1(n16383), .ip2(\pipeline/csr/from_host [1]), .op(n15838) );
  nand4_1 U17354 ( .ip1(n15841), .ip2(n15840), .ip3(n15839), .ip4(n15838), 
        .op(n15842) );
  not_ab_or_c_or_d U17355 ( .ip1(n16310), .ip2(\pipeline/csr/mtime_full [33]), 
        .ip3(n15843), .ip4(n15842), .op(n15853) );
  nand2_1 U17356 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [1]), .op(n15845)
         );
  nand2_1 U17357 ( .ip1(n16039), .ip2(\pipeline/csr/mecode [1]), .op(n15844)
         );
  nand2_1 U17358 ( .ip1(n15845), .ip2(n15844), .op(n15851) );
  nand2_1 U17359 ( .ip1(\pipeline/prv [0]), .ip2(n20964), .op(n15849) );
  nand2_1 U17360 ( .ip1(n16382), .ip2(\pipeline/csr/mtime_full [1]), .op(
        n15848) );
  nand2_1 U17361 ( .ip1(n18144), .ip2(\pipeline/csr/mie [1]), .op(n15847) );
  nand2_1 U17362 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [1]), .op(n15846)
         );
  nand4_1 U17363 ( .ip1(n15849), .ip2(n15848), .ip3(n15847), .ip4(n15846), 
        .op(n15850) );
  not_ab_or_c_or_d U17364 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [1]), 
        .ip3(n15851), .ip4(n15850), .op(n15852) );
  nand2_1 U17365 ( .ip1(n15853), .ip2(n15852), .op(n21275) );
  nand3_1 U17366 ( .ip1(n16062), .ip2(n16335), .ip3(n21275), .op(n15855) );
  nand2_1 U17367 ( .ip1(n16369), .ip2(htif_pcr_req_data[1]), .op(n15854) );
  nand2_1 U17368 ( .ip1(n15855), .ip2(n15854), .op(n16064) );
  nor2_1 U17369 ( .ip1(n15856), .ip2(n16064), .op(n22033) );
  or2_1 U17370 ( .ip1(n22033), .ip2(n15857), .op(n15861) );
  nand2_1 U17371 ( .ip1(n16413), .ip2(\pipeline/PC_WB [1]), .op(n15860) );
  nand2_1 U17372 ( .ip1(n16411), .ip2(\pipeline/csr/mbadaddr [1]), .op(n15859)
         );
  nand2_1 U17373 ( .ip1(\pipeline/alu_out_WB [1]), .ip2(n16412), .op(n15858)
         );
  nand4_1 U17374 ( .ip1(n15861), .ip2(n15860), .ip3(n15859), .ip4(n15858), 
        .op(n8699) );
  nand2_1 U17375 ( .ip1(n16368), .ip2(n20476), .op(n15891) );
  nand2_1 U17376 ( .ip1(n16369), .ip2(htif_pcr_req_data[5]), .op(n15890) );
  nand2_1 U17377 ( .ip1(n16335), .ip2(n15862), .op(n15863) );
  nand2_1 U17378 ( .ip1(n16337), .ip2(n15863), .op(n15888) );
  inv_1 U17379 ( .ip(\pipeline/csr/time_full [37]), .op(n21051) );
  nor2_1 U17380 ( .ip1(n15864), .ip2(n21051), .op(n15868) );
  nand2_1 U17381 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [5]), .op(
        n15866) );
  nand2_1 U17382 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [37]), .op(
        n15865) );
  nand2_1 U17383 ( .ip1(n15866), .ip2(n15865), .op(n15867) );
  not_ab_or_c_or_d U17384 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [5]), 
        .ip3(n15868), .ip4(n15867), .op(n15887) );
  inv_1 U17385 ( .ip(\pipeline/epc [5]), .op(n15870) );
  nor2_1 U17386 ( .ip1(n15870), .ip2(n15869), .op(n15883) );
  inv_1 U17387 ( .ip(\pipeline/csr/from_host [5]), .op(n15871) );
  nor2_1 U17388 ( .ip1(n17833), .ip2(n15871), .op(n15873) );
  inv_1 U17389 ( .ip(\pipeline/csr/instret_full [5]), .op(n17824) );
  nor2_1 U17390 ( .ip1(n16380), .ip2(n17824), .op(n15872) );
  not_ab_or_c_or_d U17391 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [5]), 
        .ip3(n15873), .ip4(n15872), .op(n15881) );
  nand2_1 U17392 ( .ip1(n20964), .ip2(\pipeline/csr/priv_stack [5]), .op(
        n15877) );
  nand2_1 U17393 ( .ip1(\pipeline/csr/mtvec [5]), .ip2(n17364), .op(n15876) );
  nand2_1 U17394 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [37]), .op(
        n15875) );
  nand2_1 U17395 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [5]), .op(n15874)
         );
  and4_1 U17396 ( .ip1(n15877), .ip2(n15876), .ip3(n15875), .ip4(n15874), .op(
        n15880) );
  nand2_1 U17397 ( .ip1(n18144), .ip2(\pipeline/csr/mie [5]), .op(n15879) );
  nand2_1 U17398 ( .ip1(n16382), .ip2(\pipeline/csr/mtime_full [5]), .op(
        n15878) );
  nand4_1 U17399 ( .ip1(n15881), .ip2(n15880), .ip3(n15879), .ip4(n15878), 
        .op(n15882) );
  not_ab_or_c_or_d U17400 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [5]), 
        .ip3(n15883), .ip4(n15882), .op(n15886) );
  nand2_1 U17401 ( .ip1(n16310), .ip2(\pipeline/csr/mtime_full [37]), .op(
        n15885) );
  nand2_1 U17402 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [5]), .op(n15884)
         );
  nand4_1 U17403 ( .ip1(n15887), .ip2(n15886), .ip3(n15885), .ip4(n15884), 
        .op(n17973) );
  nand2_1 U17404 ( .ip1(n15888), .ip2(n17973), .op(n15889) );
  nand3_1 U17405 ( .ip1(n15891), .ip2(n15890), .ip3(n15889), .op(n22145) );
  nand2_1 U17406 ( .ip1(n16410), .ip2(n22145), .op(n15895) );
  nand2_1 U17407 ( .ip1(\pipeline/csr/mbadaddr [5]), .ip2(n16411), .op(n15894)
         );
  nand2_1 U17408 ( .ip1(\pipeline/alu_out_WB [5]), .ip2(n16412), .op(n15893)
         );
  nand2_1 U17409 ( .ip1(n16413), .ip2(\pipeline/PC_WB [5]), .op(n15892) );
  nand4_1 U17410 ( .ip1(n15895), .ip2(n15894), .ip3(n15893), .ip4(n15892), 
        .op(n8695) );
  nand2_1 U17411 ( .ip1(n16368), .ip2(n15896), .op(n15923) );
  nand2_1 U17412 ( .ip1(n16369), .ip2(htif_pcr_req_data[9]), .op(n15922) );
  nand2_1 U17413 ( .ip1(n16335), .ip2(n20507), .op(n15897) );
  nand2_1 U17414 ( .ip1(n16337), .ip2(n15897), .op(n15920) );
  nand2_1 U17415 ( .ip1(ext_interrupts[1]), .ip2(n19599), .op(n15919) );
  nand2_1 U17416 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [9]), .op(n15901) );
  nand2_1 U17417 ( .ip1(n16301), .ip2(\pipeline/csr/instret_full [9]), .op(
        n15900) );
  nand2_1 U17418 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [9]), .op(n15899)
         );
  nand2_1 U17419 ( .ip1(n16383), .ip2(\pipeline/csr/from_host [9]), .op(n15898) );
  nand4_1 U17420 ( .ip1(n15901), .ip2(n15900), .ip3(n15899), .ip4(n15898), 
        .op(n15905) );
  nand2_1 U17421 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [9]), .op(n15903)
         );
  nand2_1 U17422 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [9]), .op(n15902)
         );
  nand2_1 U17423 ( .ip1(n15903), .ip2(n15902), .op(n15904) );
  not_ab_or_c_or_d U17424 ( .ip1(n16310), .ip2(\pipeline/csr/mtime_full [41]), 
        .ip3(n15905), .ip4(n15904), .op(n15918) );
  nand2_1 U17425 ( .ip1(\pipeline/csr/mie [9]), .ip2(n18144), .op(n15909) );
  nand2_1 U17426 ( .ip1(n16382), .ip2(\pipeline/csr/mtime_full [9]), .op(
        n15908) );
  nand2_1 U17427 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [9]), .op(n15907)
         );
  nand2_1 U17428 ( .ip1(\pipeline/csr/mtvec [9]), .ip2(n17364), .op(n15906) );
  nand4_1 U17429 ( .ip1(n15909), .ip2(n15908), .ip3(n15907), .ip4(n15906), 
        .op(n15915) );
  nand2_1 U17430 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [41]), .op(
        n15913) );
  nand2_1 U17431 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [9]), .op(
        n15912) );
  nand2_1 U17432 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [41]), .op(
        n15911) );
  nand2_1 U17433 ( .ip1(n16373), .ip2(\pipeline/csr/time_full [41]), .op(
        n15910) );
  nand4_1 U17434 ( .ip1(n15913), .ip2(n15912), .ip3(n15911), .ip4(n15910), 
        .op(n15914) );
  nor2_1 U17435 ( .ip1(n15915), .ip2(n15914), .op(n15917) );
  nand2_1 U17436 ( .ip1(\pipeline/epc [9]), .ip2(n17305), .op(n15916) );
  nand4_1 U17437 ( .ip1(n15919), .ip2(n15918), .ip3(n15917), .ip4(n15916), 
        .op(n19762) );
  nand2_1 U17438 ( .ip1(n15920), .ip2(n19762), .op(n15921) );
  nand3_1 U17439 ( .ip1(n15923), .ip2(n15922), .ip3(n15921), .op(n18470) );
  nand2_1 U17440 ( .ip1(n16410), .ip2(n18470), .op(n15927) );
  nand2_1 U17441 ( .ip1(\pipeline/csr/mbadaddr [9]), .ip2(n16411), .op(n15926)
         );
  nand2_1 U17442 ( .ip1(\pipeline/alu_out_WB [9]), .ip2(n16412), .op(n15925)
         );
  nand2_1 U17443 ( .ip1(n16413), .ip2(\pipeline/PC_WB [9]), .op(n15924) );
  nand4_1 U17444 ( .ip1(n15927), .ip2(n15926), .ip3(n15925), .ip4(n15924), 
        .op(n8691) );
  nand2_1 U17445 ( .ip1(n16368), .ip2(n15928), .op(n15955) );
  nand2_1 U17446 ( .ip1(n16369), .ip2(htif_pcr_req_data[7]), .op(n15954) );
  nand2_1 U17447 ( .ip1(n16335), .ip2(n20381), .op(n15929) );
  nand2_1 U17448 ( .ip1(n16337), .ip2(n15929), .op(n15952) );
  nand2_1 U17449 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [39]), .op(
        n15933) );
  nand2_1 U17450 ( .ip1(n16301), .ip2(\pipeline/csr/instret_full [7]), .op(
        n15932) );
  nand2_1 U17451 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [7]), .op(n15931)
         );
  nand2_1 U17452 ( .ip1(n16383), .ip2(\pipeline/csr/from_host [7]), .op(n15930) );
  nand4_1 U17453 ( .ip1(n15933), .ip2(n15932), .ip3(n15931), .ip4(n15930), 
        .op(n15937) );
  nand2_1 U17454 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [7]), .op(n15935)
         );
  nand2_1 U17455 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [7]), .op(n15934)
         );
  nand2_1 U17456 ( .ip1(n15935), .ip2(n15934), .op(n15936) );
  not_ab_or_c_or_d U17457 ( .ip1(n16310), .ip2(\pipeline/csr/mtime_full [39]), 
        .ip3(n15937), .ip4(n15936), .op(n15951) );
  nand2_1 U17458 ( .ip1(\pipeline/csr/mie [7]), .ip2(n18144), .op(n15941) );
  nand2_1 U17459 ( .ip1(n16382), .ip2(\pipeline/csr/mtime_full [7]), .op(
        n15940) );
  nand2_1 U17460 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [7]), .op(n15939)
         );
  nand2_1 U17461 ( .ip1(\pipeline/csr/mtvec [7]), .ip2(n17364), .op(n15938) );
  nand4_1 U17462 ( .ip1(n15941), .ip2(n15940), .ip3(n15939), .ip4(n15938), 
        .op(n15947) );
  nand2_1 U17463 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [39]), .op(
        n15945) );
  nand2_1 U17464 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [7]), .op(
        n15944) );
  nand2_1 U17465 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [7]), .op(n15943) );
  nand2_1 U17466 ( .ip1(n16373), .ip2(\pipeline/csr/time_full [39]), .op(
        n15942) );
  nand4_1 U17467 ( .ip1(n15945), .ip2(n15944), .ip3(n15943), .ip4(n15942), 
        .op(n15946) );
  nor2_1 U17468 ( .ip1(n15947), .ip2(n15946), .op(n15950) );
  nand2_1 U17469 ( .ip1(\pipeline/epc [7]), .ip2(n17305), .op(n15949) );
  nand2_1 U17470 ( .ip1(\pipeline/csr/mip[7] ), .ip2(n19599), .op(n15948) );
  nand4_1 U17471 ( .ip1(n15951), .ip2(n15950), .ip3(n15949), .ip4(n15948), 
        .op(n20390) );
  nand2_1 U17472 ( .ip1(n15952), .ip2(n20390), .op(n15953) );
  nand3_1 U17473 ( .ip1(n15955), .ip2(n15954), .ip3(n15953), .op(n19677) );
  nand2_1 U17474 ( .ip1(n16410), .ip2(n19677), .op(n15959) );
  nand2_1 U17475 ( .ip1(n16413), .ip2(\pipeline/PC_WB [7]), .op(n15958) );
  nand2_1 U17476 ( .ip1(\pipeline/csr/mbadaddr [7]), .ip2(n16411), .op(n15957)
         );
  nand2_1 U17477 ( .ip1(\pipeline/alu_out_WB [7]), .ip2(n16412), .op(n15956)
         );
  nand4_1 U17478 ( .ip1(n15959), .ip2(n15958), .ip3(n15957), .ip4(n15956), 
        .op(n8693) );
  nor2_1 U17479 ( .ip1(n15962), .ip2(n15960), .op(n15987) );
  nor2_1 U17480 ( .ip1(n15962), .ip2(n15961), .op(n15985) );
  inv_1 U17481 ( .ip(\pipeline/csr/mtime_full [38]), .op(n22153) );
  nor2_1 U17482 ( .ip1(n16338), .ip2(n22153), .op(n15983) );
  nand2_1 U17483 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [38]), .op(
        n15966) );
  nand2_1 U17484 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [6]), .op(
        n15965) );
  nand2_1 U17485 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [38]), .op(
        n15964) );
  nand2_1 U17486 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [6]), .op(n15963) );
  nand4_1 U17487 ( .ip1(n15966), .ip2(n15965), .ip3(n15964), .ip4(n15963), 
        .op(n15982) );
  nand2_1 U17488 ( .ip1(n16373), .ip2(\pipeline/csr/time_full [38]), .op(
        n15970) );
  nand2_1 U17489 ( .ip1(n16301), .ip2(\pipeline/csr/instret_full [6]), .op(
        n15969) );
  nand2_1 U17490 ( .ip1(n16383), .ip2(\pipeline/csr/from_host [6]), .op(n15968) );
  nand2_1 U17491 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [6]), .op(n15967)
         );
  nand4_1 U17492 ( .ip1(n15970), .ip2(n15969), .ip3(n15968), .ip4(n15967), 
        .op(n15981) );
  inv_1 U17493 ( .ip(\pipeline/csr/mtime_full [6]), .op(n19659) );
  nor2_1 U17494 ( .ip1(n15971), .ip2(n19659), .op(n15975) );
  nand2_1 U17495 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [6]), .op(n15973)
         );
  nand2_1 U17496 ( .ip1(\pipeline/csr/mtvec [6]), .ip2(n17364), .op(n15972) );
  nand2_1 U17497 ( .ip1(n15973), .ip2(n15972), .op(n15974) );
  not_ab_or_c_or_d U17498 ( .ip1(\pipeline/csr/mie [6]), .ip2(n18144), .ip3(
        n15975), .ip4(n15974), .op(n15979) );
  nand2_1 U17499 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [6]), .op(n15978)
         );
  nand2_1 U17500 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [6]), .op(n15977)
         );
  nand2_1 U17501 ( .ip1(\pipeline/epc [6]), .ip2(n17305), .op(n15976) );
  nand4_1 U17502 ( .ip1(n15979), .ip2(n15978), .ip3(n15977), .ip4(n15976), 
        .op(n15980) );
  nor4_1 U17503 ( .ip1(n15983), .ip2(n15982), .ip3(n15981), .ip4(n15980), .op(
        n20378) );
  nor2_1 U17504 ( .ip1(n20378), .ip2(n16401), .op(n15984) );
  nor2_1 U17505 ( .ip1(n15985), .ip2(n15984), .op(n15986) );
  or2_1 U17506 ( .ip1(n15987), .ip2(n15986), .op(n15989) );
  nand2_1 U17507 ( .ip1(n16369), .ip2(htif_pcr_req_data[6]), .op(n15988) );
  nand2_1 U17508 ( .ip1(n15989), .ip2(n15988), .op(n22364) );
  nand2_1 U17509 ( .ip1(n16410), .ip2(n22364), .op(n15993) );
  nand2_1 U17510 ( .ip1(n16411), .ip2(\pipeline/csr/mbadaddr [6]), .op(n15992)
         );
  nand2_1 U17511 ( .ip1(\pipeline/alu_out_WB [6]), .ip2(n16412), .op(n15991)
         );
  nand2_1 U17512 ( .ip1(n16413), .ip2(\pipeline/PC_WB [6]), .op(n15990) );
  nand4_1 U17513 ( .ip1(n15993), .ip2(n15992), .ip3(n15991), .ip4(n15990), 
        .op(n8694) );
  nand2_1 U17514 ( .ip1(n16310), .ip2(\pipeline/csr/mtime_full [63]), .op(
        n15997) );
  nand2_1 U17515 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [31]), .op(n15996) );
  nand2_1 U17516 ( .ip1(n16039), .ip2(\pipeline/csr/mcause[31] ), .op(n15995)
         );
  nand2_1 U17517 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [31]), .op(n15994) );
  nand4_1 U17518 ( .ip1(n15997), .ip2(n15996), .ip3(n15995), .ip4(n15994), 
        .op(n16016) );
  inv_1 U17519 ( .ip(\pipeline/csr/instret_full [31]), .op(n20956) );
  nor2_1 U17520 ( .ip1(n16380), .ip2(n20956), .op(n16002) );
  nand2_1 U17521 ( .ip1(ext_interrupts[23]), .ip2(n19599), .op(n16000) );
  nand2_1 U17522 ( .ip1(n16382), .ip2(\pipeline/csr/mtime_full [31]), .op(
        n15999) );
  nand2_1 U17523 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [31]), .op(n15998)
         );
  nand3_1 U17524 ( .ip1(n16000), .ip2(n15999), .ip3(n15998), .op(n16001) );
  not_ab_or_c_or_d U17525 ( .ip1(n16383), .ip2(\pipeline/csr/from_host [31]), 
        .ip3(n16002), .ip4(n16001), .op(n16004) );
  nand2_1 U17526 ( .ip1(\pipeline/epc [31]), .ip2(n17305), .op(n16003) );
  nand2_1 U17527 ( .ip1(n16004), .ip2(n16003), .op(n16015) );
  nand2_1 U17528 ( .ip1(\pipeline/csr/mie [31]), .ip2(n18144), .op(n16008) );
  nand2_1 U17529 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [31]), .op(n16007) );
  nand2_1 U17530 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [63]), .op(
        n16006) );
  nand2_1 U17531 ( .ip1(\pipeline/csr/mtvec [31]), .ip2(n17364), .op(n16005)
         );
  nand4_1 U17532 ( .ip1(n16008), .ip2(n16007), .ip3(n16006), .ip4(n16005), 
        .op(n16014) );
  nand2_1 U17533 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [31]), .op(
        n16012) );
  nand2_1 U17534 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [63]), .op(
        n16011) );
  nand2_1 U17535 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [31]), .op(
        n16010) );
  nand2_1 U17536 ( .ip1(n16373), .ip2(\pipeline/csr/time_full [63]), .op(
        n16009) );
  nand4_1 U17537 ( .ip1(n16012), .ip2(n16011), .ip3(n16010), .ip4(n16009), 
        .op(n16013) );
  nor4_1 U17538 ( .ip1(n16016), .ip2(n16015), .ip3(n16014), .ip4(n16013), .op(
        n21678) );
  nor2_1 U17539 ( .ip1(n14594), .ip2(n16401), .op(n16017) );
  nor2_1 U17540 ( .ip1(n16403), .ip2(n16017), .op(n16018) );
  nor2_1 U17541 ( .ip1(n21678), .ip2(n16018), .op(n16022) );
  nor3_1 U17542 ( .ip1(\pipeline/dmem_type[2] ), .ip2(n16020), .ip3(n16019), 
        .op(n16021) );
  not_ab_or_c_or_d U17543 ( .ip1(n16369), .ip2(htif_pcr_req_data[31]), .ip3(
        n16022), .ip4(n16021), .op(n22245) );
  inv_1 U17544 ( .ip(n22245), .op(n20959) );
  nand2_1 U17545 ( .ip1(n16410), .ip2(n20959), .op(n16026) );
  nand2_1 U17546 ( .ip1(n16411), .ip2(\pipeline/csr/mbadaddr [31]), .op(n16025) );
  nand2_1 U17547 ( .ip1(\pipeline/alu_out_WB [31]), .ip2(n16412), .op(n16024)
         );
  nand2_1 U17548 ( .ip1(n16413), .ip2(\pipeline/PC_WB [31]), .op(n16023) );
  nand4_1 U17549 ( .ip1(n16026), .ip2(n16025), .ip3(n16024), .ip4(n16023), 
        .op(n8669) );
  inv_1 U17550 ( .ip(n16055), .op(n16027) );
  nand2_1 U17551 ( .ip1(n20965), .ip2(n16039), .op(n16057) );
  nand3_1 U17552 ( .ip1(n16027), .ip2(n20966), .ip3(n16057), .op(n20933) );
  buf_1 U17553 ( .ip(htif_reset), .op(n21089) );
  nor2_1 U17554 ( .ip1(n21089), .ip2(n16057), .op(n21185) );
  inv_1 U17555 ( .ip(n18022), .op(n21500) );
  mux2_1 U17556 ( .ip1(n21500), .ip2(n16028), .s(\pipeline/dmem_type[2] ), 
        .op(n16052) );
  nand2_1 U17557 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [32]), .op(
        n16032) );
  nand2_1 U17558 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [0]), .op(
        n16031) );
  nand2_1 U17559 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [32]), .op(
        n16030) );
  nand2_1 U17560 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [0]), .op(n16029) );
  nand4_1 U17561 ( .ip1(n16032), .ip2(n16031), .ip3(n16030), .ip4(n16029), 
        .op(n16038) );
  nand2_1 U17562 ( .ip1(n16373), .ip2(\pipeline/csr/time_full [32]), .op(
        n16036) );
  nand2_1 U17563 ( .ip1(n16301), .ip2(\pipeline/csr/instret_full [0]), .op(
        n16035) );
  nand2_1 U17564 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [0]), .op(n16034)
         );
  nand2_1 U17565 ( .ip1(n16383), .ip2(\pipeline/csr/from_host [0]), .op(n16033) );
  nand4_1 U17566 ( .ip1(n16036), .ip2(n16035), .ip3(n16034), .ip4(n16033), 
        .op(n16037) );
  not_ab_or_c_or_d U17567 ( .ip1(n16310), .ip2(\pipeline/csr/mtime_full [32]), 
        .ip3(n16038), .ip4(n16037), .op(n16049) );
  nand2_1 U17568 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [0]), .op(n16041)
         );
  nand2_1 U17569 ( .ip1(n16039), .ip2(\pipeline/csr/mecode [0]), .op(n16040)
         );
  nand2_1 U17570 ( .ip1(n16041), .ip2(n16040), .op(n16047) );
  nand2_1 U17571 ( .ip1(n20964), .ip2(\pipeline/csr/priv_stack_0 ), .op(n16045) );
  nand2_1 U17572 ( .ip1(n16382), .ip2(\pipeline/csr/mtime_full [0]), .op(
        n16044) );
  nand2_1 U17573 ( .ip1(n18144), .ip2(\pipeline/csr/mie [0]), .op(n16043) );
  nand2_1 U17574 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [0]), .op(n16042)
         );
  nand4_1 U17575 ( .ip1(n16045), .ip2(n16044), .ip3(n16043), .ip4(n16042), 
        .op(n16046) );
  not_ab_or_c_or_d U17576 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [0]), 
        .ip3(n16047), .ip4(n16046), .op(n16048) );
  nand2_1 U17577 ( .ip1(n16049), .ip2(n16048), .op(n21527) );
  nand3_1 U17578 ( .ip1(n16052), .ip2(n16335), .ip3(n21527), .op(n16051) );
  nand2_1 U17579 ( .ip1(n16369), .ip2(htif_pcr_req_data[0]), .op(n16050) );
  and2_1 U17580 ( .ip1(n16051), .ip2(n16050), .op(n16075) );
  inv_1 U17581 ( .ip(n16052), .op(n16072) );
  nand2_1 U17582 ( .ip1(n17949), .ip2(n16072), .op(n16053) );
  nand2_1 U17583 ( .ip1(n16075), .ip2(n16053), .op(n22377) );
  nand2_1 U17584 ( .ip1(n21185), .ip2(n22377), .op(n16061) );
  nor2_1 U17585 ( .ip1(n21089), .ip2(n20972), .op(n16054) );
  nand3_1 U17586 ( .ip1(n16055), .ip2(n16054), .ip3(n16057), .op(n16066) );
  nor2_1 U17587 ( .ip1(n16056), .ip2(n16066), .op(n21187) );
  nand2_1 U17588 ( .ip1(n21187), .ip2(\pipeline/ctrl/prev_ex_code_WB [0]), 
        .op(n16060) );
  nor2_1 U17589 ( .ip1(n21089), .ip2(n10364), .op(n16058) );
  nand2_1 U17590 ( .ip1(n16058), .ip2(n16057), .op(n21125) );
  inv_1 U17591 ( .ip(n21125), .op(n21186) );
  nand2_1 U17592 ( .ip1(n21186), .ip2(\pipeline/csr/mecode [0]), .op(n16059)
         );
  nand4_1 U17593 ( .ip1(n20933), .ip2(n16061), .ip3(n16060), .ip4(n16059), 
        .op(n8735) );
  inv_1 U17594 ( .ip(n17949), .op(n16063) );
  nor2_1 U17595 ( .ip1(n16063), .ip2(n16062), .op(n16065) );
  nor2_1 U17596 ( .ip1(n16065), .ip2(n16064), .op(n22261) );
  inv_1 U17597 ( .ip(n22261), .op(n22129) );
  nand2_1 U17598 ( .ip1(n21185), .ip2(n22129), .op(n16071) );
  nand2_1 U17599 ( .ip1(n21187), .ip2(\pipeline/ctrl/prev_ex_code_WB [1]), 
        .op(n16070) );
  nand2_1 U17600 ( .ip1(n21186), .ip2(\pipeline/csr/mecode [1]), .op(n16069)
         );
  nor2_1 U17601 ( .ip1(\pipeline/ctrl/had_ex_WB ), .ip2(n16066), .op(n21128)
         );
  inv_1 U17602 ( .ip(\pipeline/ctrl/wr_reg_unkilled_WB ), .op(n16067) );
  nand2_1 U17603 ( .ip1(n21128), .ip2(n16067), .op(n16068) );
  nand4_1 U17604 ( .ip1(n16071), .ip2(n16070), .ip3(n16069), .ip4(n16068), 
        .op(n8734) );
  nand2_1 U17605 ( .ip1(n16073), .ip2(n16072), .op(n16074) );
  nand2_1 U17606 ( .ip1(n16075), .ip2(n16074), .op(n16076) );
  nand2_1 U17607 ( .ip1(n16410), .ip2(n16076), .op(n16080) );
  nand2_1 U17608 ( .ip1(n16413), .ip2(\pipeline/PC_WB [0]), .op(n16079) );
  nand2_1 U17609 ( .ip1(n16411), .ip2(\pipeline/csr/mbadaddr [0]), .op(n16078)
         );
  nand2_1 U17610 ( .ip1(\pipeline/alu_out_WB [0]), .ip2(n16412), .op(n16077)
         );
  nand4_1 U17611 ( .ip1(n16080), .ip2(n16079), .ip3(n16078), .ip4(n16077), 
        .op(n8700) );
  nand2_1 U17612 ( .ip1(n16368), .ip2(n14593), .op(n16107) );
  nand2_1 U17613 ( .ip1(n16369), .ip2(htif_pcr_req_data[16]), .op(n16106) );
  nand2_1 U17614 ( .ip1(n16335), .ip2(n18148), .op(n16081) );
  nand2_1 U17615 ( .ip1(n16337), .ip2(n16081), .op(n16104) );
  nand2_1 U17616 ( .ip1(ext_interrupts[8]), .ip2(n19599), .op(n16103) );
  nand2_1 U17617 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [48]), .op(
        n16085) );
  nand2_1 U17618 ( .ip1(n16301), .ip2(\pipeline/csr/instret_full [16]), .op(
        n16084) );
  nand2_1 U17619 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [16]), .op(n16083)
         );
  nand2_1 U17620 ( .ip1(n16383), .ip2(\pipeline/csr/from_host [16]), .op(
        n16082) );
  nand4_1 U17621 ( .ip1(n16085), .ip2(n16084), .ip3(n16083), .ip4(n16082), 
        .op(n16089) );
  nand2_1 U17622 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [16]), .op(n16087) );
  nand2_1 U17623 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [16]), .op(n16086) );
  nand2_1 U17624 ( .ip1(n16087), .ip2(n16086), .op(n16088) );
  not_ab_or_c_or_d U17625 ( .ip1(n16310), .ip2(\pipeline/csr/mtime_full [48]), 
        .ip3(n16089), .ip4(n16088), .op(n16102) );
  nand2_1 U17626 ( .ip1(\pipeline/csr/mie [16]), .ip2(n18144), .op(n16093) );
  nand2_1 U17627 ( .ip1(n16382), .ip2(\pipeline/csr/mtime_full [16]), .op(
        n16092) );
  nand2_1 U17628 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [16]), .op(n16091) );
  nand2_1 U17629 ( .ip1(\pipeline/csr/mtvec [16]), .ip2(n17364), .op(n16090)
         );
  nand4_1 U17630 ( .ip1(n16093), .ip2(n16092), .ip3(n16091), .ip4(n16090), 
        .op(n16099) );
  nand2_1 U17631 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [48]), .op(
        n16097) );
  nand2_1 U17632 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [16]), .op(
        n16096) );
  nand2_1 U17633 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [16]), .op(
        n16095) );
  nand2_1 U17634 ( .ip1(n16373), .ip2(\pipeline/csr/time_full [48]), .op(
        n16094) );
  nand4_1 U17635 ( .ip1(n16097), .ip2(n16096), .ip3(n16095), .ip4(n16094), 
        .op(n16098) );
  nor2_1 U17636 ( .ip1(n16099), .ip2(n16098), .op(n16101) );
  nand2_1 U17637 ( .ip1(\pipeline/epc [16]), .ip2(n17305), .op(n16100) );
  nand4_1 U17638 ( .ip1(n16103), .ip2(n16102), .ip3(n16101), .ip4(n16100), 
        .op(n19956) );
  nand2_1 U17639 ( .ip1(n16104), .ip2(n19956), .op(n16105) );
  nand3_1 U17640 ( .ip1(n16107), .ip2(n16106), .ip3(n16105), .op(n19951) );
  nand2_1 U17641 ( .ip1(n16410), .ip2(n19951), .op(n16111) );
  nand2_1 U17642 ( .ip1(\pipeline/csr/mbadaddr [16]), .ip2(n16411), .op(n16110) );
  nand2_1 U17643 ( .ip1(\pipeline/alu_out_WB [16]), .ip2(n16412), .op(n16109)
         );
  nand2_1 U17644 ( .ip1(n16413), .ip2(\pipeline/PC_WB [16]), .op(n16108) );
  nand4_1 U17645 ( .ip1(n16111), .ip2(n16110), .ip3(n16109), .ip4(n16108), 
        .op(n8684) );
  nand2_1 U17646 ( .ip1(n16368), .ip2(n20611), .op(n16139) );
  nand2_1 U17647 ( .ip1(n16369), .ip2(htif_pcr_req_data[24]), .op(n16138) );
  nand2_1 U17648 ( .ip1(n16335), .ip2(n16112), .op(n16113) );
  nand2_1 U17649 ( .ip1(n16337), .ip2(n16113), .op(n16136) );
  nand2_1 U17650 ( .ip1(ext_interrupts[16]), .ip2(n19599), .op(n16135) );
  nand2_1 U17651 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [56]), .op(
        n16117) );
  nand2_1 U17652 ( .ip1(n16301), .ip2(\pipeline/csr/instret_full [24]), .op(
        n16116) );
  nand2_1 U17653 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [24]), .op(n16115)
         );
  nand2_1 U17654 ( .ip1(n16383), .ip2(\pipeline/csr/from_host [24]), .op(
        n16114) );
  nand4_1 U17655 ( .ip1(n16117), .ip2(n16116), .ip3(n16115), .ip4(n16114), 
        .op(n16121) );
  nand2_1 U17656 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [24]), .op(n16119) );
  nand2_1 U17657 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [24]), .op(n16118) );
  nand2_1 U17658 ( .ip1(n16119), .ip2(n16118), .op(n16120) );
  not_ab_or_c_or_d U17659 ( .ip1(n16310), .ip2(\pipeline/csr/mtime_full [56]), 
        .ip3(n16121), .ip4(n16120), .op(n16134) );
  nand2_1 U17660 ( .ip1(\pipeline/csr/mie [24]), .ip2(n18144), .op(n16125) );
  nand2_1 U17661 ( .ip1(n16382), .ip2(\pipeline/csr/mtime_full [24]), .op(
        n16124) );
  nand2_1 U17662 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [24]), .op(n16123) );
  nand2_1 U17663 ( .ip1(\pipeline/csr/mtvec [24]), .ip2(n17364), .op(n16122)
         );
  nand4_1 U17664 ( .ip1(n16125), .ip2(n16124), .ip3(n16123), .ip4(n16122), 
        .op(n16131) );
  nand2_1 U17665 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [56]), .op(
        n16129) );
  nand2_1 U17666 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [24]), .op(
        n16128) );
  nand2_1 U17667 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [24]), .op(
        n16127) );
  nand2_1 U17668 ( .ip1(n16373), .ip2(\pipeline/csr/time_full [56]), .op(
        n16126) );
  nand4_1 U17669 ( .ip1(n16129), .ip2(n16128), .ip3(n16127), .ip4(n16126), 
        .op(n16130) );
  nor2_1 U17670 ( .ip1(n16131), .ip2(n16130), .op(n16133) );
  nand2_1 U17671 ( .ip1(\pipeline/epc [24]), .ip2(n17305), .op(n16132) );
  nand4_1 U17672 ( .ip1(n16135), .ip2(n16134), .ip3(n16133), .ip4(n16132), 
        .op(n21985) );
  nand2_1 U17673 ( .ip1(n16136), .ip2(n21985), .op(n16137) );
  nand3_1 U17674 ( .ip1(n16139), .ip2(n16138), .ip3(n16137), .op(n18794) );
  nand2_1 U17675 ( .ip1(n16410), .ip2(n18794), .op(n16143) );
  nand2_1 U17676 ( .ip1(\pipeline/csr/mbadaddr [24]), .ip2(n16411), .op(n16142) );
  nand2_1 U17677 ( .ip1(\pipeline/alu_out_WB [24]), .ip2(n16412), .op(n16141)
         );
  nand2_1 U17678 ( .ip1(n16413), .ip2(\pipeline/PC_WB [24]), .op(n16140) );
  nand4_1 U17679 ( .ip1(n16143), .ip2(n16142), .ip3(n16141), .ip4(n16140), 
        .op(n8676) );
  nand2_1 U17680 ( .ip1(n16368), .ip2(n20646), .op(n16170) );
  and2_1 U17681 ( .ip1(n16369), .ip2(htif_pcr_req_data[28]), .op(n16168) );
  and2_1 U17682 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [28]), .op(n16164)
         );
  inv_1 U17683 ( .ip(\pipeline/csr/mtime_full [60]), .op(n22231) );
  nor2_1 U17684 ( .ip1(n16338), .ip2(n22231), .op(n16163) );
  nand2_1 U17685 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [28]), .op(
        n16147) );
  nand2_1 U17686 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [60]), .op(
        n16146) );
  nand2_1 U17687 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [28]), .op(
        n16145) );
  nand2_1 U17688 ( .ip1(n16373), .ip2(\pipeline/csr/time_full [60]), .op(
        n16144) );
  nand4_1 U17689 ( .ip1(n16147), .ip2(n16146), .ip3(n16145), .ip4(n16144), 
        .op(n16162) );
  inv_1 U17690 ( .ip(\pipeline/csr/instret_full [28]), .op(n19287) );
  nor2_1 U17691 ( .ip1(n16380), .ip2(n19287), .op(n16152) );
  nand2_1 U17692 ( .ip1(ext_interrupts[20]), .ip2(n19599), .op(n16150) );
  nand2_1 U17693 ( .ip1(n16382), .ip2(\pipeline/csr/mtime_full [28]), .op(
        n16149) );
  nand2_1 U17694 ( .ip1(n16383), .ip2(\pipeline/csr/from_host [28]), .op(
        n16148) );
  nand3_1 U17695 ( .ip1(n16150), .ip2(n16149), .ip3(n16148), .op(n16151) );
  not_ab_or_c_or_d U17696 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [28]), 
        .ip3(n16152), .ip4(n16151), .op(n16160) );
  nand2_1 U17697 ( .ip1(\pipeline/csr/mie [28]), .ip2(n18144), .op(n16156) );
  nand2_1 U17698 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [28]), .op(n16155) );
  nand2_1 U17699 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [60]), .op(
        n16154) );
  nand2_1 U17700 ( .ip1(\pipeline/csr/mtvec [28]), .ip2(n17364), .op(n16153)
         );
  and4_1 U17701 ( .ip1(n16156), .ip2(n16155), .ip3(n16154), .ip4(n16153), .op(
        n16159) );
  nand2_1 U17702 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [28]), .op(n16158) );
  nand2_1 U17703 ( .ip1(\pipeline/epc [28]), .ip2(n17305), .op(n16157) );
  nand4_1 U17704 ( .ip1(n16160), .ip2(n16159), .ip3(n16158), .ip4(n16157), 
        .op(n16161) );
  nor4_1 U17705 ( .ip1(n16164), .ip2(n16163), .ip3(n16162), .ip4(n16161), .op(
        n19299) );
  nor2_1 U17706 ( .ip1(n20646), .ip2(n16401), .op(n16165) );
  nor2_1 U17707 ( .ip1(n16165), .ip2(n16403), .op(n16166) );
  nor2_1 U17708 ( .ip1(n19299), .ip2(n16166), .op(n16167) );
  nor2_1 U17709 ( .ip1(n16168), .ip2(n16167), .op(n16169) );
  and2_1 U17710 ( .ip1(n16170), .ip2(n16169), .op(n22229) );
  inv_1 U17711 ( .ip(n22229), .op(n22281) );
  nand2_1 U17712 ( .ip1(n16410), .ip2(n22281), .op(n16174) );
  nand2_1 U17713 ( .ip1(\pipeline/csr/mbadaddr [28]), .ip2(n16411), .op(n16173) );
  nand2_1 U17714 ( .ip1(\pipeline/alu_out_WB [28]), .ip2(n16412), .op(n16172)
         );
  nand2_1 U17715 ( .ip1(n16413), .ip2(\pipeline/PC_WB [28]), .op(n16171) );
  nand4_1 U17716 ( .ip1(n16174), .ip2(n16173), .ip3(n16172), .ip4(n16171), 
        .op(n8672) );
  nand2_1 U17717 ( .ip1(n16368), .ip2(n21645), .op(n16199) );
  and2_1 U17718 ( .ip1(n16369), .ip2(htif_pcr_req_data[30]), .op(n16197) );
  nand2_1 U17719 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [30]), .op(
        n16178) );
  nand2_1 U17720 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [62]), .op(
        n16177) );
  nand2_1 U17721 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [30]), .op(
        n16176) );
  nand2_1 U17722 ( .ip1(n16373), .ip2(\pipeline/csr/time_full [62]), .op(
        n16175) );
  and4_1 U17723 ( .ip1(n16178), .ip2(n16177), .ip3(n16176), .ip4(n16175), .op(
        n16195) );
  inv_1 U17724 ( .ip(\pipeline/csr/instret_full [30]), .op(n19006) );
  nor2_1 U17725 ( .ip1(n16380), .ip2(n19006), .op(n16183) );
  nand2_1 U17726 ( .ip1(ext_interrupts[22]), .ip2(n19599), .op(n16181) );
  nand2_1 U17727 ( .ip1(n16382), .ip2(\pipeline/csr/mtime_full [30]), .op(
        n16180) );
  nand2_1 U17728 ( .ip1(n16383), .ip2(\pipeline/csr/from_host [30]), .op(
        n16179) );
  nand3_1 U17729 ( .ip1(n16181), .ip2(n16180), .ip3(n16179), .op(n16182) );
  not_ab_or_c_or_d U17730 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [30]), 
        .ip3(n16183), .ip4(n16182), .op(n16191) );
  nand2_1 U17731 ( .ip1(\pipeline/csr/mie [30]), .ip2(n18144), .op(n16187) );
  nand2_1 U17732 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [30]), .op(n16186) );
  nand2_1 U17733 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [62]), .op(
        n16185) );
  nand2_1 U17734 ( .ip1(\pipeline/csr/mtvec [30]), .ip2(n17364), .op(n16184)
         );
  and4_1 U17735 ( .ip1(n16187), .ip2(n16186), .ip3(n16185), .ip4(n16184), .op(
        n16190) );
  nand2_1 U17736 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [30]), .op(n16189) );
  nand2_1 U17737 ( .ip1(\pipeline/epc [30]), .ip2(n17305), .op(n16188) );
  and4_1 U17738 ( .ip1(n16191), .ip2(n16190), .ip3(n16189), .ip4(n16188), .op(
        n16194) );
  nand2_1 U17739 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [30]), .op(n16193) );
  nand2_1 U17740 ( .ip1(n16310), .ip2(\pipeline/csr/mtime_full [62]), .op(
        n16192) );
  and4_1 U17741 ( .ip1(n16195), .ip2(n16194), .ip3(n16193), .ip4(n16192), .op(
        n19011) );
  not_ab_or_c_or_d U17742 ( .ip1(n17765), .ip2(n21645), .ip3(n19011), .ip4(
        n16401), .op(n16196) );
  nor2_1 U17743 ( .ip1(n16197), .ip2(n16196), .op(n16198) );
  and2_1 U17744 ( .ip1(n16199), .ip2(n16198), .op(n22258) );
  inv_1 U17745 ( .ip(n22258), .op(n22313) );
  nand2_1 U17746 ( .ip1(n16410), .ip2(n22313), .op(n16203) );
  nand2_1 U17747 ( .ip1(\pipeline/csr/mbadaddr [30]), .ip2(n16411), .op(n16202) );
  nand2_1 U17748 ( .ip1(\pipeline/alu_out_WB [30]), .ip2(n16412), .op(n16201)
         );
  nand2_1 U17749 ( .ip1(n16413), .ip2(\pipeline/PC_WB [30]), .op(n16200) );
  nand4_1 U17750 ( .ip1(n16203), .ip2(n16202), .ip3(n16201), .ip4(n16200), 
        .op(n8670) );
  nand2_1 U17751 ( .ip1(n16368), .ip2(n16226), .op(n16232) );
  and2_1 U17752 ( .ip1(n16369), .ip2(htif_pcr_req_data[11]), .op(n16230) );
  nand2_1 U17753 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [43]), .op(
        n16207) );
  nand2_1 U17754 ( .ip1(n16301), .ip2(\pipeline/csr/instret_full [11]), .op(
        n16206) );
  nand2_1 U17755 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [11]), .op(n16205)
         );
  nand2_1 U17756 ( .ip1(n16383), .ip2(\pipeline/csr/from_host [11]), .op(
        n16204) );
  nand4_1 U17757 ( .ip1(n16207), .ip2(n16206), .ip3(n16205), .ip4(n16204), 
        .op(n16211) );
  nand2_1 U17758 ( .ip1(\pipeline/epc [11]), .ip2(n17305), .op(n16209) );
  nand2_1 U17759 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [11]), .op(n16208) );
  nand2_1 U17760 ( .ip1(n16209), .ip2(n16208), .op(n16210) );
  not_ab_or_c_or_d U17761 ( .ip1(n16310), .ip2(\pipeline/csr/mtime_full [43]), 
        .ip3(n16211), .ip4(n16210), .op(n16225) );
  nand2_1 U17762 ( .ip1(\pipeline/csr/mie [11]), .ip2(n18144), .op(n16215) );
  nand2_1 U17763 ( .ip1(n16382), .ip2(\pipeline/csr/mtime_full [11]), .op(
        n16214) );
  nand2_1 U17764 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [11]), .op(n16213) );
  nand2_1 U17765 ( .ip1(\pipeline/csr/mtvec [11]), .ip2(n17364), .op(n16212)
         );
  nand4_1 U17766 ( .ip1(n16215), .ip2(n16214), .ip3(n16213), .ip4(n16212), 
        .op(n16221) );
  nand2_1 U17767 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [43]), .op(
        n16219) );
  nand2_1 U17768 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [11]), .op(
        n16218) );
  nand2_1 U17769 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [11]), .op(
        n16217) );
  nand2_1 U17770 ( .ip1(n16373), .ip2(\pipeline/csr/time_full [43]), .op(
        n16216) );
  nand4_1 U17771 ( .ip1(n16219), .ip2(n16218), .ip3(n16217), .ip4(n16216), 
        .op(n16220) );
  nor2_1 U17772 ( .ip1(n16221), .ip2(n16220), .op(n16224) );
  nand2_1 U17773 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [11]), .op(n16223) );
  nand2_1 U17774 ( .ip1(ext_interrupts[3]), .ip2(n19599), .op(n16222) );
  and4_1 U17775 ( .ip1(n16225), .ip2(n16224), .ip3(n16223), .ip4(n16222), .op(
        n20201) );
  nor2_1 U17776 ( .ip1(n16226), .ip2(n16401), .op(n16227) );
  nor2_1 U17777 ( .ip1(n16227), .ip2(n16403), .op(n16228) );
  nor2_1 U17778 ( .ip1(n20201), .ip2(n16228), .op(n16229) );
  nor2_1 U17779 ( .ip1(n16230), .ip2(n16229), .op(n16231) );
  and2_1 U17780 ( .ip1(n16232), .ip2(n16231), .op(n20196) );
  inv_1 U17781 ( .ip(n20196), .op(n22156) );
  nand2_1 U17782 ( .ip1(n16410), .ip2(n22156), .op(n16236) );
  nand2_1 U17783 ( .ip1(\pipeline/csr/mbadaddr [11]), .ip2(n16411), .op(n16235) );
  nand2_1 U17784 ( .ip1(\pipeline/alu_out_WB [11]), .ip2(n16412), .op(n16234)
         );
  nand2_1 U17785 ( .ip1(n16413), .ip2(\pipeline/PC_WB [11]), .op(n16233) );
  nand4_1 U17786 ( .ip1(n16236), .ip2(n16235), .ip3(n16234), .ip4(n16233), 
        .op(n8689) );
  nand2_1 U17787 ( .ip1(n16368), .ip2(n16237), .op(n16265) );
  nand2_1 U17788 ( .ip1(n16369), .ip2(htif_pcr_req_data[27]), .op(n16264) );
  nand2_1 U17789 ( .ip1(n16335), .ip2(n16238), .op(n16239) );
  nand2_1 U17790 ( .ip1(n16337), .ip2(n16239), .op(n16262) );
  nand2_1 U17791 ( .ip1(ext_interrupts[19]), .ip2(n19599), .op(n16261) );
  nand2_1 U17792 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [27]), .op(
        n16243) );
  nand2_1 U17793 ( .ip1(n16301), .ip2(\pipeline/csr/instret_full [27]), .op(
        n16242) );
  nand2_1 U17794 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [27]), .op(n16241)
         );
  nand2_1 U17795 ( .ip1(n16383), .ip2(\pipeline/csr/from_host [27]), .op(
        n16240) );
  nand4_1 U17796 ( .ip1(n16243), .ip2(n16242), .ip3(n16241), .ip4(n16240), 
        .op(n16247) );
  nand2_1 U17797 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [27]), .op(n16245) );
  nand2_1 U17798 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [27]), .op(n16244) );
  nand2_1 U17799 ( .ip1(n16245), .ip2(n16244), .op(n16246) );
  not_ab_or_c_or_d U17800 ( .ip1(n16310), .ip2(\pipeline/csr/mtime_full [59]), 
        .ip3(n16247), .ip4(n16246), .op(n16260) );
  nand2_1 U17801 ( .ip1(\pipeline/csr/mie [27]), .ip2(n18144), .op(n16251) );
  nand2_1 U17802 ( .ip1(n16382), .ip2(\pipeline/csr/mtime_full [27]), .op(
        n16250) );
  nand2_1 U17803 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [27]), .op(n16249) );
  nand2_1 U17804 ( .ip1(\pipeline/csr/mtvec [27]), .ip2(n17364), .op(n16248)
         );
  nand4_1 U17805 ( .ip1(n16251), .ip2(n16250), .ip3(n16249), .ip4(n16248), 
        .op(n16257) );
  nand2_1 U17806 ( .ip1(n16373), .ip2(\pipeline/csr/time_full [59]), .op(
        n16255) );
  nand2_1 U17807 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [59]), .op(
        n16254) );
  nand2_1 U17808 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [27]), .op(
        n16253) );
  nand2_1 U17809 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [59]), .op(
        n16252) );
  nand4_1 U17810 ( .ip1(n16255), .ip2(n16254), .ip3(n16253), .ip4(n16252), 
        .op(n16256) );
  nor2_1 U17811 ( .ip1(n16257), .ip2(n16256), .op(n16259) );
  nand2_1 U17812 ( .ip1(\pipeline/epc [27]), .ip2(n17305), .op(n16258) );
  nand4_1 U17813 ( .ip1(n16261), .ip2(n16260), .ip3(n16259), .ip4(n16258), 
        .op(n20163) );
  nand2_1 U17814 ( .ip1(n16262), .ip2(n20163), .op(n16263) );
  nand3_1 U17815 ( .ip1(n16265), .ip2(n16264), .ip3(n16263), .op(n19243) );
  nand2_1 U17816 ( .ip1(n16410), .ip2(n19243), .op(n16269) );
  nand2_1 U17817 ( .ip1(n16413), .ip2(\pipeline/PC_WB [27]), .op(n16268) );
  nand2_1 U17818 ( .ip1(\pipeline/csr/mbadaddr [27]), .ip2(n16411), .op(n16267) );
  nand2_1 U17819 ( .ip1(\pipeline/alu_out_WB [27]), .ip2(n16412), .op(n16266)
         );
  nand4_1 U17820 ( .ip1(n16269), .ip2(n16268), .ip3(n16267), .ip4(n16266), 
        .op(n8673) );
  nand2_1 U17821 ( .ip1(n16368), .ip2(n20650), .op(n16296) );
  nand2_1 U17822 ( .ip1(n16369), .ip2(htif_pcr_req_data[29]), .op(n16295) );
  nand2_1 U17823 ( .ip1(n16335), .ip2(n21622), .op(n16270) );
  nand2_1 U17824 ( .ip1(n16337), .ip2(n16270), .op(n16293) );
  nand2_1 U17825 ( .ip1(ext_interrupts[21]), .ip2(n19599), .op(n16292) );
  nand2_1 U17826 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [61]), .op(
        n16274) );
  nand2_1 U17827 ( .ip1(n16301), .ip2(\pipeline/csr/instret_full [29]), .op(
        n16273) );
  nand2_1 U17828 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [29]), .op(n16272)
         );
  nand2_1 U17829 ( .ip1(n16383), .ip2(\pipeline/csr/from_host [29]), .op(
        n16271) );
  nand4_1 U17830 ( .ip1(n16274), .ip2(n16273), .ip3(n16272), .ip4(n16271), 
        .op(n16278) );
  nand2_1 U17831 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [29]), .op(n16276) );
  nand2_1 U17832 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [29]), .op(n16275) );
  nand2_1 U17833 ( .ip1(n16276), .ip2(n16275), .op(n16277) );
  not_ab_or_c_or_d U17834 ( .ip1(n16310), .ip2(\pipeline/csr/mtime_full [61]), 
        .ip3(n16278), .ip4(n16277), .op(n16291) );
  nand2_1 U17835 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [29]), .op(n16282) );
  nand2_1 U17836 ( .ip1(n16382), .ip2(\pipeline/csr/mtime_full [29]), .op(
        n16281) );
  nand2_1 U17837 ( .ip1(\pipeline/csr/mie [29]), .ip2(n18144), .op(n16280) );
  nand2_1 U17838 ( .ip1(\pipeline/csr/mtvec [29]), .ip2(n17364), .op(n16279)
         );
  nand4_1 U17839 ( .ip1(n16282), .ip2(n16281), .ip3(n16280), .ip4(n16279), 
        .op(n16288) );
  nand2_1 U17840 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [61]), .op(
        n16286) );
  nand2_1 U17841 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [29]), .op(
        n16285) );
  nand2_1 U17842 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [29]), .op(
        n16284) );
  nand2_1 U17843 ( .ip1(n16373), .ip2(\pipeline/csr/time_full [61]), .op(
        n16283) );
  nand4_1 U17844 ( .ip1(n16286), .ip2(n16285), .ip3(n16284), .ip4(n16283), 
        .op(n16287) );
  nor2_1 U17845 ( .ip1(n16288), .ip2(n16287), .op(n16290) );
  nand2_1 U17846 ( .ip1(\pipeline/epc [29]), .ip2(n17305), .op(n16289) );
  nand4_1 U17847 ( .ip1(n16292), .ip2(n16291), .ip3(n16290), .ip4(n16289), 
        .op(n20688) );
  nand2_1 U17848 ( .ip1(n16293), .ip2(n20688), .op(n16294) );
  nand3_1 U17849 ( .ip1(n16296), .ip2(n16295), .ip3(n16294), .op(n22234) );
  nand2_1 U17850 ( .ip1(n16410), .ip2(n22234), .op(n16300) );
  nand2_1 U17851 ( .ip1(\pipeline/csr/mbadaddr [29]), .ip2(n16411), .op(n16299) );
  nand2_1 U17852 ( .ip1(\pipeline/alu_out_WB [29]), .ip2(n16412), .op(n16298)
         );
  nand2_1 U17853 ( .ip1(n16413), .ip2(\pipeline/PC_WB [29]), .op(n16297) );
  nand4_1 U17854 ( .ip1(n16300), .ip2(n16299), .ip3(n16298), .ip4(n16297), 
        .op(n8671) );
  nand2_1 U17855 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [42]), .op(
        n16305) );
  nand2_1 U17856 ( .ip1(n16301), .ip2(\pipeline/csr/instret_full [10]), .op(
        n16304) );
  nand2_1 U17857 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [10]), .op(n16303)
         );
  nand2_1 U17858 ( .ip1(n16383), .ip2(\pipeline/csr/from_host [10]), .op(
        n16302) );
  nand4_1 U17859 ( .ip1(n16305), .ip2(n16304), .ip3(n16303), .ip4(n16302), 
        .op(n16309) );
  nand2_1 U17860 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [10]), .op(n16307) );
  nand2_1 U17861 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [10]), .op(n16306) );
  nand2_1 U17862 ( .ip1(n16307), .ip2(n16306), .op(n16308) );
  not_ab_or_c_or_d U17863 ( .ip1(n16310), .ip2(\pipeline/csr/mtime_full [42]), 
        .ip3(n16309), .ip4(n16308), .op(n16324) );
  nand2_1 U17864 ( .ip1(\pipeline/csr/mie [10]), .ip2(n18144), .op(n16314) );
  nand2_1 U17865 ( .ip1(n16382), .ip2(\pipeline/csr/mtime_full [10]), .op(
        n16313) );
  nand2_1 U17866 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [10]), .op(n16312) );
  nand2_1 U17867 ( .ip1(\pipeline/csr/mtvec [10]), .ip2(n17364), .op(n16311)
         );
  nand4_1 U17868 ( .ip1(n16314), .ip2(n16313), .ip3(n16312), .ip4(n16311), 
        .op(n16320) );
  nand2_1 U17869 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [42]), .op(
        n16318) );
  nand2_1 U17870 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [10]), .op(
        n16317) );
  nand2_1 U17871 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [10]), .op(
        n16316) );
  nand2_1 U17872 ( .ip1(n16373), .ip2(\pipeline/csr/time_full [42]), .op(
        n16315) );
  nand4_1 U17873 ( .ip1(n16318), .ip2(n16317), .ip3(n16316), .ip4(n16315), 
        .op(n16319) );
  nor2_1 U17874 ( .ip1(n16320), .ip2(n16319), .op(n16323) );
  nand2_1 U17875 ( .ip1(\pipeline/epc [10]), .ip2(n17305), .op(n16322) );
  nand2_1 U17876 ( .ip1(ext_interrupts[2]), .ip2(n19599), .op(n16321) );
  and4_1 U17877 ( .ip1(n16324), .ip2(n16323), .ip3(n16322), .ip4(n16321), .op(
        n19833) );
  nor2_1 U17878 ( .ip1(n14601), .ip2(n16401), .op(n16325) );
  nor2_1 U17879 ( .ip1(n16325), .ip2(n16403), .op(n16326) );
  nor2_1 U17880 ( .ip1(n19833), .ip2(n16326), .op(n16328) );
  and2_1 U17881 ( .ip1(n16369), .ip2(htif_pcr_req_data[10]), .op(n16327) );
  not_ab_or_c_or_d U17882 ( .ip1(n16368), .ip2(n14601), .ip3(n16328), .ip4(
        n16327), .op(n19805) );
  inv_1 U17883 ( .ip(n19805), .op(n19828) );
  nand2_1 U17884 ( .ip1(n16410), .ip2(n19828), .op(n16332) );
  nand2_1 U17885 ( .ip1(\pipeline/csr/mbadaddr [10]), .ip2(n16411), .op(n16331) );
  nand2_1 U17886 ( .ip1(\pipeline/alu_out_WB [10]), .ip2(n16412), .op(n16330)
         );
  nand2_1 U17887 ( .ip1(n16413), .ip2(\pipeline/PC_WB [10]), .op(n16329) );
  nand4_1 U17888 ( .ip1(n16332), .ip2(n16331), .ip3(n16330), .ip4(n16329), 
        .op(n8690) );
  nand2_1 U17889 ( .ip1(n16368), .ip2(n16333), .op(n16363) );
  nand2_1 U17890 ( .ip1(n16369), .ip2(htif_pcr_req_data[26]), .op(n16362) );
  nand2_1 U17891 ( .ip1(n16335), .ip2(n16334), .op(n16336) );
  nand2_1 U17892 ( .ip1(n16337), .ip2(n16336), .op(n16360) );
  inv_1 U17893 ( .ip(\pipeline/csr/mtime_full [58]), .op(n22226) );
  nor2_1 U17894 ( .ip1(n16338), .ip2(n22226), .op(n16344) );
  nand2_1 U17895 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [26]), .op(
        n16342) );
  nand2_1 U17896 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [58]), .op(
        n16341) );
  nand2_1 U17897 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [26]), .op(
        n16340) );
  nand2_1 U17898 ( .ip1(n16373), .ip2(\pipeline/csr/time_full [58]), .op(
        n16339) );
  nand4_1 U17899 ( .ip1(n16342), .ip2(n16341), .ip3(n16340), .ip4(n16339), 
        .op(n16343) );
  not_ab_or_c_or_d U17900 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [26]), 
        .ip3(n16344), .ip4(n16343), .op(n16359) );
  inv_1 U17901 ( .ip(\pipeline/csr/instret_full [26]), .op(n19125) );
  nor2_1 U17902 ( .ip1(n16380), .ip2(n19125), .op(n16355) );
  and2_1 U17903 ( .ip1(n22096), .ip2(\pipeline/csr/to_host [26]), .op(n16354)
         );
  nand2_1 U17904 ( .ip1(ext_interrupts[18]), .ip2(n19599), .op(n16347) );
  nand2_1 U17905 ( .ip1(n16382), .ip2(\pipeline/csr/mtime_full [26]), .op(
        n16346) );
  nand2_1 U17906 ( .ip1(n16383), .ip2(\pipeline/csr/from_host [26]), .op(
        n16345) );
  nand3_1 U17907 ( .ip1(n16347), .ip2(n16346), .ip3(n16345), .op(n16353) );
  nand2_1 U17908 ( .ip1(\pipeline/csr/mie [26]), .ip2(n18144), .op(n16351) );
  nand2_1 U17909 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [26]), .op(n16350) );
  nand2_1 U17910 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [58]), .op(
        n16349) );
  nand2_1 U17911 ( .ip1(\pipeline/csr/mtvec [26]), .ip2(n17364), .op(n16348)
         );
  nand4_1 U17912 ( .ip1(n16351), .ip2(n16350), .ip3(n16349), .ip4(n16348), 
        .op(n16352) );
  nor4_1 U17913 ( .ip1(n16355), .ip2(n16354), .ip3(n16353), .ip4(n16352), .op(
        n16358) );
  nand2_1 U17914 ( .ip1(\pipeline/epc [26]), .ip2(n17305), .op(n16357) );
  nand2_1 U17915 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [26]), .op(n16356) );
  nand4_1 U17916 ( .ip1(n16359), .ip2(n16358), .ip3(n16357), .ip4(n16356), 
        .op(n20315) );
  nand2_1 U17917 ( .ip1(n16360), .ip2(n20315), .op(n16361) );
  nand3_1 U17918 ( .ip1(n16363), .ip2(n16362), .ip3(n16361), .op(n22222) );
  nand2_1 U17919 ( .ip1(n16410), .ip2(n22222), .op(n16367) );
  nand2_1 U17920 ( .ip1(\pipeline/csr/mbadaddr [26]), .ip2(n16411), .op(n16366) );
  nand2_1 U17921 ( .ip1(\pipeline/alu_out_WB [26]), .ip2(n16412), .op(n16365)
         );
  nand2_1 U17922 ( .ip1(n16413), .ip2(\pipeline/PC_WB [26]), .op(n16364) );
  nand4_1 U17923 ( .ip1(n16367), .ip2(n16366), .ip3(n16365), .ip4(n16364), 
        .op(n8674) );
  nand2_1 U17924 ( .ip1(n16368), .ip2(n16402), .op(n16409) );
  and2_1 U17925 ( .ip1(n16369), .ip2(htif_pcr_req_data[12]), .op(n16407) );
  inv_1 U17926 ( .ip(\pipeline/csr/mtime_full [44]), .op(n22163) );
  nor2_1 U17927 ( .ip1(n16338), .ip2(n22163), .op(n16379) );
  nand2_1 U17928 ( .ip1(n16370), .ip2(\pipeline/csr/cycle_full [12]), .op(
        n16377) );
  nand2_1 U17929 ( .ip1(n16371), .ip2(\pipeline/csr/instret_full [44]), .op(
        n16376) );
  nand2_1 U17930 ( .ip1(n16372), .ip2(\pipeline/csr/time_full [12]), .op(
        n16375) );
  nand2_1 U17931 ( .ip1(n16373), .ip2(\pipeline/csr/time_full [44]), .op(
        n16374) );
  nand4_1 U17932 ( .ip1(n16377), .ip2(n16376), .ip3(n16375), .ip4(n16374), 
        .op(n16378) );
  not_ab_or_c_or_d U17933 ( .ip1(n17828), .ip2(\pipeline/csr/mscratch [12]), 
        .ip3(n16379), .ip4(n16378), .op(n16400) );
  inv_1 U17934 ( .ip(\pipeline/csr/instret_full [12]), .op(n20781) );
  nor2_1 U17935 ( .ip1(n16380), .ip2(n20781), .op(n16395) );
  inv_1 U17936 ( .ip(\pipeline/csr/to_host [12]), .op(n16381) );
  nor2_1 U17937 ( .ip1(n17843), .ip2(n16381), .op(n16394) );
  nand2_1 U17938 ( .ip1(ext_interrupts[4]), .ip2(n19599), .op(n16386) );
  nand2_1 U17939 ( .ip1(n16382), .ip2(\pipeline/csr/mtime_full [12]), .op(
        n16385) );
  nand2_1 U17940 ( .ip1(n16383), .ip2(\pipeline/csr/from_host [12]), .op(
        n16384) );
  nand3_1 U17941 ( .ip1(n16386), .ip2(n16385), .ip3(n16384), .op(n16393) );
  nand2_1 U17942 ( .ip1(\pipeline/csr/mie [12]), .ip2(n18144), .op(n16391) );
  nand2_1 U17943 ( .ip1(n17812), .ip2(\pipeline/csr/mtimecmp [12]), .op(n16390) );
  nand2_1 U17944 ( .ip1(n16387), .ip2(\pipeline/csr/cycle_full [44]), .op(
        n16389) );
  nand2_1 U17945 ( .ip1(\pipeline/csr/mtvec [12]), .ip2(n17364), .op(n16388)
         );
  nand4_1 U17946 ( .ip1(n16391), .ip2(n16390), .ip3(n16389), .ip4(n16388), 
        .op(n16392) );
  nor4_1 U17947 ( .ip1(n16395), .ip2(n16394), .ip3(n16393), .ip4(n16392), .op(
        n16399) );
  nand2_1 U17948 ( .ip1(\pipeline/epc [12]), .ip2(n17305), .op(n16398) );
  nand2_1 U17949 ( .ip1(n16396), .ip2(\pipeline/csr/mbadaddr [12]), .op(n16397) );
  and4_1 U17950 ( .ip1(n16400), .ip2(n16399), .ip3(n16398), .ip4(n16397), .op(
        n20794) );
  nor2_1 U17951 ( .ip1(n16402), .ip2(n16401), .op(n16404) );
  nor2_1 U17952 ( .ip1(n16404), .ip2(n16403), .op(n16405) );
  nor2_1 U17953 ( .ip1(n20794), .ip2(n16405), .op(n16406) );
  nor2_1 U17954 ( .ip1(n16407), .ip2(n16406), .op(n16408) );
  nand2_1 U17955 ( .ip1(n16409), .ip2(n16408), .op(n20788) );
  nand2_1 U17956 ( .ip1(n16410), .ip2(n20788), .op(n16417) );
  nand2_1 U17957 ( .ip1(\pipeline/csr/mbadaddr [12]), .ip2(n16411), .op(n16416) );
  nand2_1 U17958 ( .ip1(\pipeline/alu_out_WB [12]), .ip2(n16412), .op(n16415)
         );
  nand2_1 U17959 ( .ip1(n16413), .ip2(\pipeline/PC_WB [12]), .op(n16414) );
  nand4_1 U17960 ( .ip1(n16417), .ip2(n16416), .ip3(n16415), .ip4(n16414), 
        .op(n8688) );
  xor2_1 U17961 ( .ip1(n16418), .ip2(n16913), .op(n16419) );
  nor2_1 U17962 ( .ip1(n16419), .ip2(n16845), .op(n16574) );
  inv_1 U17963 ( .ip(n16574), .op(n16565) );
  nand2_1 U17964 ( .ip1(n16419), .ip2(n16845), .op(n16567) );
  nand2_1 U17965 ( .ip1(n16565), .ip2(n16567), .op(n16476) );
  xor2_1 U17966 ( .ip1(n19432), .ip2(n20855), .op(n16437) );
  nand2_1 U17967 ( .ip1(n16437), .ip2(n19433), .op(n19415) );
  inv_1 U17968 ( .ip(n19415), .op(n16564) );
  xor2_1 U17969 ( .ip1(n16913), .ip2(n17142), .op(n16420) );
  nand2_1 U17970 ( .ip1(n16420), .ip2(n12138), .op(n17128) );
  nor2_1 U17971 ( .ip1(n16420), .ip2(n12138), .op(n16434) );
  inv_1 U17972 ( .ip(n16434), .op(n17129) );
  xor2_1 U17973 ( .ip1(n20222), .ip2(n20855), .op(n16433) );
  nand2_1 U17974 ( .ip1(n16433), .ip2(n20221), .op(n20207) );
  inv_1 U17975 ( .ip(n20207), .op(n17132) );
  nand2_1 U17976 ( .ip1(n17129), .ip2(n17132), .op(n16421) );
  nand2_1 U17977 ( .ip1(n17128), .ip2(n16421), .op(n16436) );
  xor2_1 U17978 ( .ip1(n20728), .ip2(n16913), .op(n16422) );
  nand2_1 U17979 ( .ip1(n16422), .ip2(n13627), .op(n20708) );
  inv_1 U17980 ( .ip(n20708), .op(n16425) );
  nor2_1 U17981 ( .ip1(n16422), .ip2(n16838), .op(n16427) );
  xor2_1 U17982 ( .ip1(n16690), .ip2(n20855), .op(n16426) );
  nand2_1 U17983 ( .ip1(n16426), .ip2(n16423), .op(n20710) );
  nor2_1 U17984 ( .ip1(n16427), .ip2(n20710), .op(n16424) );
  nor2_1 U17985 ( .ip1(n16425), .ip2(n16424), .op(n16432) );
  nor2_1 U17986 ( .ip1(n16426), .ip2(n16423), .op(n20711) );
  inv_1 U17987 ( .ip(n20711), .op(n20715) );
  inv_1 U17988 ( .ip(n16427), .op(n20709) );
  nand2_1 U17989 ( .ip1(n20715), .ip2(n20709), .op(n16441) );
  xor2_1 U17990 ( .ip1(n16972), .ip2(n16913), .op(n16428) );
  nand2_1 U17991 ( .ip1(n16428), .ip2(n16973), .op(n16962) );
  inv_1 U17992 ( .ip(n16962), .op(n16430) );
  nor2_1 U17993 ( .ip1(n16428), .ip2(n16973), .op(n16440) );
  xor2_1 U17994 ( .ip1(n17457), .ip2(n20855), .op(n16439) );
  nand2_1 U17995 ( .ip1(n16439), .ip2(n17456), .op(n17468) );
  nor2_1 U17996 ( .ip1(n16440), .ip2(n17468), .op(n16429) );
  nor2_1 U17997 ( .ip1(n16430), .ip2(n16429), .op(n20712) );
  or2_1 U17998 ( .ip1(n16441), .ip2(n20712), .op(n16431) );
  nand2_1 U17999 ( .ip1(n16432), .ip2(n16431), .op(n17130) );
  nor2_1 U18000 ( .ip1(n16433), .ip2(n20221), .op(n17133) );
  nor2_1 U18001 ( .ip1(n16434), .ip2(n17133), .op(n16442) );
  and2_1 U18002 ( .ip1(n17130), .ip2(n16442), .op(n16435) );
  nor2_1 U18003 ( .ip1(n16436), .ip2(n16435), .op(n19419) );
  nor2_1 U18004 ( .ip1(n16437), .ip2(n19433), .op(n16573) );
  nor2_1 U18005 ( .ip1(n19419), .ip2(n16573), .op(n16438) );
  nor2_1 U18006 ( .ip1(n16564), .ip2(n16438), .op(n16474) );
  nor2_1 U18007 ( .ip1(n16439), .ip2(n17456), .op(n16964) );
  inv_1 U18008 ( .ip(n16964), .op(n17469) );
  inv_1 U18009 ( .ip(n16440), .op(n16963) );
  nand2_1 U18010 ( .ip1(n17469), .ip2(n16963), .op(n16665) );
  nor2_1 U18011 ( .ip1(n16665), .ip2(n16441), .op(n20209) );
  nand2_1 U18012 ( .ip1(n20209), .ip2(n16442), .op(n16578) );
  inv_1 U18013 ( .ip(n16578), .op(n19417) );
  inv_1 U18014 ( .ip(n16573), .op(n19416) );
  nand2_1 U18015 ( .ip1(n19417), .ip2(n19416), .op(n16472) );
  nand2_1 U18016 ( .ip1(n16443), .ip2(n10185), .op(n17191) );
  xor2_1 U18017 ( .ip1(n16776), .ip2(n16913), .op(n16459) );
  nand2_1 U18018 ( .ip1(n16459), .ip2(n17492), .op(n16750) );
  inv_1 U18019 ( .ip(n16750), .op(n17194) );
  nor2_1 U18020 ( .ip1(n16443), .ip2(n10185), .op(n16460) );
  inv_1 U18021 ( .ip(n16460), .op(n17192) );
  nand2_1 U18022 ( .ip1(n17194), .ip2(n17192), .op(n16444) );
  nand2_1 U18023 ( .ip1(n17191), .ip2(n16444), .op(n17567) );
  xor2_1 U18024 ( .ip1(n12596), .ip2(n16913), .op(n16452) );
  nor2_1 U18025 ( .ip1(n16452), .ip2(n13698), .op(n16454) );
  inv_1 U18026 ( .ip(n16454), .op(n16789) );
  inv_1 U18027 ( .ip(n16791), .op(n16988) );
  nand2_1 U18028 ( .ip1(n16789), .ip2(n16988), .op(n16451) );
  xor2_1 U18029 ( .ip1(n16913), .ip2(n17584), .op(n16447) );
  nor2_1 U18030 ( .ip1(n16445), .ip2(n16447), .op(n17561) );
  xor2_1 U18031 ( .ip1(n17040), .ip2(n16913), .op(n16448) );
  nor2_1 U18032 ( .ip1(n16448), .ip2(n12932), .op(n17020) );
  nor2_1 U18033 ( .ip1(n17561), .ip2(n17020), .op(n16990) );
  inv_1 U18034 ( .ip(n16990), .op(n16991) );
  nor2_1 U18035 ( .ip1(n16451), .ip2(n16991), .op(n16461) );
  nand2_1 U18036 ( .ip1(n16447), .ip2(n10187), .op(n17562) );
  nor2_1 U18037 ( .ip1(n17020), .ip2(n17562), .op(n16450) );
  nand2_1 U18038 ( .ip1(n16448), .ip2(n12932), .op(n17021) );
  inv_1 U18039 ( .ip(n17021), .op(n16449) );
  nor2_1 U18040 ( .ip1(n16450), .ip2(n16449), .op(n16995) );
  nor2_1 U18041 ( .ip1(n16451), .ip2(n16995), .op(n16458) );
  nand2_1 U18042 ( .ip1(n16452), .ip2(n13698), .op(n16788) );
  inv_1 U18043 ( .ip(n16788), .op(n16456) );
  nand2_1 U18044 ( .ip1(n16453), .ip2(n13022), .op(n16987) );
  nor2_1 U18045 ( .ip1(n16454), .ip2(n16987), .op(n16455) );
  or2_1 U18046 ( .ip1(n16456), .ip2(n16455), .op(n16457) );
  not_ab_or_c_or_d U18047 ( .ip1(n17567), .ip2(n16461), .ip3(n16458), .ip4(
        n16457), .op(n16471) );
  nor2_1 U18048 ( .ip1(n16459), .ip2(n17492), .op(n17193) );
  nor2_1 U18049 ( .ip1(n17193), .ip2(n16460), .op(n16794) );
  nand2_1 U18050 ( .ip1(n16461), .ip2(n16794), .op(n16469) );
  xor2_1 U18051 ( .ip1(n10198), .ip2(n16913), .op(n16462) );
  nand2_1 U18052 ( .ip1(n16462), .ip2(n10184), .op(n16707) );
  xor2_1 U18053 ( .ip1(n16913), .ip2(n16732), .op(n16465) );
  nand2_1 U18054 ( .ip1(n16465), .ip2(n17479), .op(n17504) );
  nor2_1 U18055 ( .ip1(n16462), .ip2(n10184), .op(n16706) );
  or2_1 U18056 ( .ip1(n17504), .ip2(n16706), .op(n16463) );
  nand2_1 U18057 ( .ip1(n16707), .ip2(n16463), .op(n16468) );
  xor2_1 U18058 ( .ip1(n16487), .ip2(n20855), .op(n21575) );
  or2_1 U18059 ( .ip1(n13524), .ip2(n16913), .op(n21574) );
  nand2_1 U18060 ( .ip1(n21575), .ip2(n21574), .op(n16464) );
  nand2_1 U18061 ( .ip1(n13524), .ip2(n16913), .op(n21573) );
  nand2_1 U18062 ( .ip1(n16464), .ip2(n21573), .op(n17503) );
  nor2_1 U18063 ( .ip1(n16465), .ip2(n17479), .op(n16704) );
  nor2_1 U18064 ( .ip1(n16706), .ip2(n16704), .op(n16466) );
  nor2_1 U18065 ( .ip1(n16468), .ip2(n16467), .op(n17565) );
  or2_1 U18066 ( .ip1(n16469), .ip2(n17565), .op(n16470) );
  nand2_1 U18067 ( .ip1(n16471), .ip2(n16470), .op(n20210) );
  inv_1 U18068 ( .ip(n20210), .op(n20717) );
  or2_1 U18069 ( .ip1(n16472), .ip2(n20717), .op(n16473) );
  nand2_1 U18070 ( .ip1(n16474), .ip2(n16473), .op(n16475) );
  xnor2_1 U18071 ( .ip1(n16476), .ip2(n16475), .op(n16486) );
  nor3_1 U18072 ( .ip1(\pipeline/dmem_type[2] ), .ip2(n16478), .ip3(n16477), 
        .op(n16482) );
  nor2_1 U18073 ( .ip1(n16480), .ip2(n16479), .op(n16481) );
  nor2_1 U18074 ( .ip1(n16482), .ip2(n16481), .op(n16484) );
  nor2_1 U18075 ( .ip1(n16484), .ip2(n16483), .op(n21530) );
  nor2_1 U18076 ( .ip1(n21530), .ip2(n16485), .op(n21577) );
  nand2_1 U18077 ( .ip1(n16486), .ip2(n21577), .op(n16541) );
  nor2_1 U18078 ( .ip1(n21530), .ip2(n16913), .op(n16524) );
  nand2_1 U18079 ( .ip1(n13894), .ip2(n16524), .op(n16501) );
  or2_1 U18080 ( .ip1(n16501), .ip2(n17199), .op(n20724) );
  nor2_1 U18081 ( .ip1(n13881), .ip2(n20724), .op(n16522) );
  and2_1 U18082 ( .ip1(n16522), .ip2(n10198), .op(n18374) );
  inv_1 U18083 ( .ip(n17480), .op(n17097) );
  and2_1 U18084 ( .ip1(n17097), .ip2(n21552), .op(n20892) );
  nand2_1 U18085 ( .ip1(n20892), .ip2(n10195), .op(n16489) );
  inv_1 U18086 ( .ip(n16507), .op(n21532) );
  inv_1 U18087 ( .ip(n21532), .op(n18927) );
  nand2_1 U18088 ( .ip1(n13540), .ip2(n18927), .op(n16488) );
  nand2_1 U18089 ( .ip1(n16489), .ip2(n16488), .op(n16491) );
  mux2_1 U18090 ( .ip1(n10184), .ip2(n17479), .s(n21552), .op(n17035) );
  nor2_1 U18091 ( .ip1(n17097), .ip2(n17035), .op(n16490) );
  nor2_1 U18092 ( .ip1(n16491), .ip2(n16490), .op(n17235) );
  inv_1 U18093 ( .ip(n16496), .op(n16493) );
  inv_1 U18094 ( .ip(n16524), .op(n16492) );
  nor2_1 U18095 ( .ip1(n16493), .ip2(n16492), .op(n20911) );
  or2_1 U18096 ( .ip1(n21555), .ip2(n16495), .op(n16505) );
  inv_1 U18097 ( .ip(n21530), .op(n16497) );
  nand3_1 U18098 ( .ip1(n16496), .ip2(n16913), .ip3(n16497), .op(n20907) );
  inv_1 U18099 ( .ip(n20907), .op(n21557) );
  nand2_1 U18100 ( .ip1(n13868), .ip2(n16498), .op(n16500) );
  nand3_1 U18101 ( .ip1(n16525), .ip2(n16913), .ip3(n16497), .op(n21551) );
  nor3_1 U18102 ( .ip1(n16498), .ip2(n21551), .ip3(n13868), .op(n16499) );
  nand2_1 U18103 ( .ip1(n13894), .ip2(n16913), .op(n16523) );
  inv_1 U18104 ( .ip(n16523), .op(n20902) );
  and2_1 U18105 ( .ip1(n17199), .ip2(n20902), .op(n20239) );
  nand2_1 U18106 ( .ip1(n20239), .ip2(n20856), .op(n20735) );
  inv_1 U18107 ( .ip(n20735), .op(n19066) );
  not_ab_or_c_or_d U18108 ( .ip1(n21557), .ip2(n16500), .ip3(n16499), .ip4(
        n19066), .op(n16504) );
  or2_1 U18109 ( .ip1(n10198), .ip2(n13525), .op(n17443) );
  inv_1 U18110 ( .ip(n21552), .op(n21553) );
  nand2_1 U18111 ( .ip1(n13524), .ip2(n21553), .op(n21534) );
  nor2_1 U18112 ( .ip1(n17443), .ip2(n21534), .op(n21563) );
  inv_1 U18113 ( .ip(n16501), .op(n16502) );
  nand2_1 U18114 ( .ip1(n17199), .ip2(n16502), .op(n20883) );
  nor2_1 U18115 ( .ip1(n16776), .ip2(n20883), .op(n17547) );
  nand2_1 U18116 ( .ip1(n21563), .ip2(n17547), .op(n16503) );
  nand3_1 U18117 ( .ip1(n16505), .ip2(n16504), .ip3(n16503), .op(n16515) );
  nand2_1 U18118 ( .ip1(n21553), .ip2(n17480), .op(n17268) );
  inv_1 U18119 ( .ip(n17268), .op(n21536) );
  nand2_1 U18120 ( .ip1(n21536), .ip2(n12138), .op(n16509) );
  nand2_1 U18121 ( .ip1(n18927), .ip2(n16845), .op(n16508) );
  nand2_1 U18122 ( .ip1(n16509), .ip2(n16508), .op(n16513) );
  nand2_1 U18123 ( .ip1(n20892), .ip2(n16846), .op(n16511) );
  nand2_1 U18124 ( .ip1(n21552), .ip2(n16732), .op(n17267) );
  inv_1 U18125 ( .ip(n17267), .op(n19056) );
  nand2_1 U18126 ( .ip1(n19056), .ip2(n20221), .op(n16510) );
  nand2_1 U18127 ( .ip1(n16511), .ip2(n16510), .op(n16512) );
  nor2_1 U18128 ( .ip1(n16513), .ip2(n16512), .op(n19060) );
  nor2_1 U18129 ( .ip1(n16776), .ip2(n20724), .op(n21562) );
  inv_1 U18130 ( .ip(n10198), .op(n17575) );
  and2_1 U18131 ( .ip1(n21562), .ip2(n17575), .op(n17541) );
  inv_1 U18132 ( .ip(n17541), .op(n17275) );
  nor2_1 U18133 ( .ip1(n19060), .ip2(n17275), .op(n16514) );
  not_ab_or_c_or_d U18134 ( .ip1(n18374), .ip2(n17235), .ip3(n16515), .ip4(
        n16514), .op(n16540) );
  and2_1 U18135 ( .ip1(n21562), .ip2(n10198), .op(n17529) );
  nand2_1 U18136 ( .ip1(n21536), .ip2(n13877), .op(n16804) );
  nand2_1 U18137 ( .ip1(n10189), .ip2(n18927), .op(n16516) );
  nand2_1 U18138 ( .ip1(n16804), .ip2(n16516), .op(n16518) );
  nand2_1 U18139 ( .ip1(n20892), .ip2(n13552), .op(n16733) );
  or2_1 U18140 ( .ip1(n17456), .ip2(n17267), .op(n16737) );
  nand2_1 U18141 ( .ip1(n16733), .ip2(n16737), .op(n16517) );
  nor2_1 U18142 ( .ip1(n16518), .ip2(n16517), .op(n19046) );
  nor2_1 U18143 ( .ip1(n10187), .ip2(n17267), .op(n16520) );
  nor2_1 U18144 ( .ip1(n12932), .ip2(n17268), .op(n16519) );
  nor2_1 U18145 ( .ip1(n16520), .ip2(n16519), .op(n16521) );
  inv_1 U18146 ( .ip(n13698), .op(n16811) );
  nand2_1 U18147 ( .ip1(n16811), .ip2(n18927), .op(n16805) );
  nand2_1 U18148 ( .ip1(n20892), .ip2(n10193), .op(n16738) );
  nand3_1 U18149 ( .ip1(n16521), .ip2(n16805), .ip3(n16738), .op(n19050) );
  and2_1 U18150 ( .ip1(n16522), .ip2(n17575), .op(n18367) );
  inv_1 U18151 ( .ip(n18367), .op(n16873) );
  nor2_1 U18152 ( .ip1(n19050), .ip2(n16873), .op(n16532) );
  or2_1 U18153 ( .ip1(n16523), .ip2(n17199), .op(n17558) );
  nand2_1 U18154 ( .ip1(n16525), .ip2(n16524), .op(n16672) );
  or2_1 U18155 ( .ip1(n16672), .ip2(n17199), .op(n19186) );
  nand2_1 U18156 ( .ip1(n17558), .ip2(n19186), .op(n21572) );
  and2_1 U18157 ( .ip1(n21572), .ip2(n13881), .op(n20736) );
  inv_1 U18158 ( .ip(n20736), .op(n17498) );
  nand2_1 U18159 ( .ip1(n16732), .ip2(n10198), .op(n17237) );
  inv_1 U18160 ( .ip(n10849), .op(n18737) );
  mux2_1 U18161 ( .ip1(n18737), .ip2(n18738), .s(n21552), .op(n17222) );
  nor2_1 U18162 ( .ip1(n17237), .ip2(n17222), .op(n16530) );
  nand2_1 U18163 ( .ip1(n17480), .ip2(n17575), .op(n17223) );
  mux2_1 U18164 ( .ip1(n16684), .ip2(n10188), .s(n21552), .op(n17208) );
  nor2_1 U18165 ( .ip1(n17223), .ip2(n17208), .op(n16529) );
  mux2_1 U18166 ( .ip1(n16845), .ip2(n16627), .s(n21552), .op(n17207) );
  nor2_1 U18167 ( .ip1(n17443), .ip2(n17207), .op(n16528) );
  nor2_1 U18168 ( .ip1(n17575), .ip2(n16732), .op(n17543) );
  inv_1 U18169 ( .ip(n17543), .op(n17227) );
  inv_1 U18170 ( .ip(n10192), .op(n17530) );
  mux2_1 U18171 ( .ip1(n17270), .ip2(n17530), .s(n21552), .op(n17225) );
  nor2_1 U18172 ( .ip1(n17227), .ip2(n17225), .op(n16527) );
  or4_1 U18173 ( .ip1(n16530), .ip2(n16529), .ip3(n16528), .ip4(n16527), .op(
        n21564) );
  nor2_1 U18174 ( .ip1(n17498), .ip2(n21564), .op(n16531) );
  not_ab_or_c_or_d U18175 ( .ip1(n17529), .ip2(n19046), .ip3(n16532), .ip4(
        n16531), .op(n16539) );
  inv_1 U18176 ( .ip(n16533), .op(n19199) );
  mux2_1 U18177 ( .ip1(n19051), .ip2(n19199), .s(n21552), .op(n17224) );
  nor2_1 U18178 ( .ip1(n17223), .ip2(n17224), .op(n21548) );
  mux2_1 U18179 ( .ip1(n10186), .ip2(n16914), .s(n21552), .op(n17226) );
  nor2_1 U18180 ( .ip1(n17443), .ip2(n17226), .op(n21547) );
  inv_1 U18181 ( .ip(n10191), .op(n20891) );
  nand2_1 U18182 ( .ip1(n20892), .ip2(n10191), .op(n16535) );
  nand2_1 U18183 ( .ip1(n10180), .ip2(n18927), .op(n16534) );
  nand2_1 U18184 ( .ip1(n16535), .ip2(n16534), .op(n16537) );
  mux2_1 U18185 ( .ip1(n17073), .ip2(n20856), .s(n21552), .op(n17121) );
  nor2_1 U18186 ( .ip1(n17097), .ip2(n17121), .op(n16536) );
  nor2_1 U18187 ( .ip1(n16537), .ip2(n16536), .op(n20733) );
  nor2_1 U18188 ( .ip1(n17575), .ip2(n20733), .op(n21545) );
  nor3_1 U18189 ( .ip1(n21548), .ip2(n21547), .ip3(n21545), .op(n18729) );
  and2_1 U18190 ( .ip1(n21572), .ip2(n16776), .op(n21549) );
  nand2_1 U18191 ( .ip1(n18729), .ip2(n21549), .op(n16538) );
  xor2_1 U18192 ( .ip1(n16594), .ip2(n20855), .op(n16542) );
  nor2_1 U18193 ( .ip1(n16542), .ip2(n18738), .op(n16924) );
  inv_1 U18194 ( .ip(n16924), .op(n16543) );
  nand2_1 U18195 ( .ip1(n16542), .ip2(n18738), .op(n16919) );
  nand2_1 U18196 ( .ip1(n16543), .ip2(n16919), .op(n16585) );
  xor2_1 U18197 ( .ip1(n17173), .ip2(n20855), .op(n16544) );
  nand2_1 U18198 ( .ip1(n16544), .ip2(n18737), .op(n17159) );
  inv_1 U18199 ( .ip(n17159), .op(n16547) );
  nor2_1 U18200 ( .ip1(n16544), .ip2(n18737), .op(n16548) );
  xor2_1 U18201 ( .ip1(n16545), .ip2(n20855), .op(n16549) );
  nand2_1 U18202 ( .ip1(n16549), .ip2(n17530), .op(n17515) );
  nor2_1 U18203 ( .ip1(n16548), .ip2(n17515), .op(n16546) );
  nor2_1 U18204 ( .ip1(n16547), .ip2(n16546), .op(n16917) );
  inv_1 U18205 ( .ip(n16548), .op(n17160) );
  nor2_1 U18206 ( .ip1(n16549), .ip2(n17530), .op(n17161) );
  inv_1 U18207 ( .ip(n17161), .op(n17516) );
  nand2_1 U18208 ( .ip1(n17160), .ip2(n17516), .op(n16925) );
  xor2_1 U18209 ( .ip1(n16550), .ip2(n20855), .op(n16551) );
  nand2_1 U18210 ( .ip1(n16551), .ip2(n17270), .op(n17243) );
  inv_1 U18211 ( .ip(n17243), .op(n16554) );
  nor2_1 U18212 ( .ip1(n16551), .ip2(n17270), .op(n16555) );
  xor2_1 U18213 ( .ip1(n16552), .ip2(n20855), .op(n16556) );
  nand2_1 U18214 ( .ip1(n16556), .ip2(n10188), .op(n17245) );
  nor2_1 U18215 ( .ip1(n16555), .ip2(n17245), .op(n16553) );
  nor2_1 U18216 ( .ip1(n16554), .ip2(n16553), .op(n16563) );
  inv_1 U18217 ( .ip(n16555), .op(n17244) );
  nor2_1 U18218 ( .ip1(n16556), .ip2(n10188), .op(n17246) );
  inv_1 U18219 ( .ip(n17246), .op(n17250) );
  nand2_1 U18220 ( .ip1(n17244), .ip2(n17250), .op(n16570) );
  xor2_1 U18221 ( .ip1(n16557), .ip2(n16913), .op(n16558) );
  nand2_1 U18222 ( .ip1(n16558), .ip2(n16854), .op(n16824) );
  inv_1 U18223 ( .ip(n16824), .op(n16561) );
  nor2_1 U18224 ( .ip1(n16558), .ip2(n16684), .op(n16568) );
  xor2_1 U18225 ( .ip1(n16913), .ip2(n16559), .op(n16569) );
  nand2_1 U18226 ( .ip1(n16569), .ip2(n16627), .op(n16827) );
  nor2_1 U18227 ( .ip1(n16568), .ip2(n16827), .op(n16560) );
  nor2_1 U18228 ( .ip1(n16561), .ip2(n16560), .op(n17247) );
  or2_1 U18229 ( .ip1(n16570), .ip2(n17247), .op(n16562) );
  nand2_1 U18230 ( .ip1(n16563), .ip2(n16562), .op(n16572) );
  nand2_1 U18231 ( .ip1(n16565), .ip2(n16564), .op(n16566) );
  nand2_1 U18232 ( .ip1(n16567), .ip2(n16566), .op(n16880) );
  inv_1 U18233 ( .ip(n16568), .op(n16825) );
  nor2_1 U18234 ( .ip1(n16569), .ip2(n16627), .op(n16828) );
  inv_1 U18235 ( .ip(n16828), .op(n16617) );
  nand2_1 U18236 ( .ip1(n16825), .ip2(n16617), .op(n16882) );
  nor2_1 U18237 ( .ip1(n16570), .ip2(n16882), .op(n16575) );
  and2_1 U18238 ( .ip1(n16880), .ip2(n16575), .op(n16571) );
  nor2_1 U18239 ( .ip1(n16572), .ip2(n16571), .op(n16577) );
  nor2_1 U18240 ( .ip1(n16574), .ip2(n16573), .op(n16619) );
  nand2_1 U18241 ( .ip1(n16575), .ip2(n16619), .op(n16579) );
  or2_1 U18242 ( .ip1(n16579), .ip2(n19419), .op(n16576) );
  nand2_1 U18243 ( .ip1(n16577), .ip2(n16576), .op(n16582) );
  nor2_1 U18244 ( .ip1(n16579), .ip2(n16578), .op(n16580) );
  and2_1 U18245 ( .ip1(n20210), .ip2(n16580), .op(n16581) );
  or2_1 U18246 ( .ip1(n16582), .ip2(n16581), .op(n20878) );
  inv_1 U18247 ( .ip(n20878), .op(n19177) );
  or2_1 U18248 ( .ip1(n16925), .ip2(n19177), .op(n16583) );
  nand2_1 U18249 ( .ip1(n16917), .ip2(n16583), .op(n16584) );
  xnor2_1 U18250 ( .ip1(n16585), .ip2(n16584), .op(n16586) );
  nand2_1 U18251 ( .ip1(n16586), .ip2(n21577), .op(n16616) );
  nand2_1 U18252 ( .ip1(n21536), .ip2(n16627), .op(n16687) );
  nand2_1 U18253 ( .ip1(n18927), .ip2(n10188), .op(n16678) );
  nand2_1 U18254 ( .ip1(n20892), .ip2(n16684), .op(n16660) );
  nand2_1 U18255 ( .ip1(n19056), .ip2(n16626), .op(n16587) );
  nand2_1 U18256 ( .ip1(n21536), .ip2(n17530), .op(n16679) );
  nand2_1 U18257 ( .ip1(n18927), .ip2(n18738), .op(n16612) );
  nand2_1 U18258 ( .ip1(n20892), .ip2(n18737), .op(n16657) );
  nand2_1 U18259 ( .ip1(n19056), .ip2(n17270), .op(n16659) );
  and4_1 U18260 ( .ip1(n16679), .ip2(n16612), .ip3(n16657), .ip4(n16659), .op(
        n20897) );
  nor2_1 U18261 ( .ip1(n17275), .ip2(n20897), .op(n16605) );
  nor2_1 U18262 ( .ip1(n13552), .ip2(n21532), .op(n16589) );
  inv_1 U18263 ( .ip(n20892), .op(n17269) );
  nor2_1 U18264 ( .ip1(n13877), .ip2(n17269), .op(n16588) );
  nor2_1 U18265 ( .ip1(n17267), .ip2(n16811), .op(n17486) );
  nor2_1 U18266 ( .ip1(n10206), .ip2(n17268), .op(n16763) );
  inv_1 U18267 ( .ip(n19422), .op(n16894) );
  nand2_1 U18268 ( .ip1(n21536), .ip2(n20221), .op(n16592) );
  nand2_1 U18269 ( .ip1(n18927), .ip2(n19433), .op(n16686) );
  nand2_1 U18270 ( .ip1(n20892), .ip2(n12138), .op(n16591) );
  nand2_1 U18271 ( .ip1(n19056), .ip2(n16838), .op(n16590) );
  inv_1 U18272 ( .ip(n19426), .op(n19194) );
  nor2_1 U18273 ( .ip1(n16873), .ip2(n19194), .op(n16603) );
  nor3_1 U18274 ( .ip1(n16593), .ip2(n21551), .ip3(n13654), .op(n16597) );
  nor2_1 U18275 ( .ip1(n16594), .ip2(n18738), .op(n16595) );
  nor2_1 U18276 ( .ip1(n20907), .ip2(n16595), .op(n16596) );
  not_ab_or_c_or_d U18277 ( .ip1(n20911), .ip2(n16598), .ip3(n16597), .ip4(
        n16596), .op(n16601) );
  nand3_1 U18278 ( .ip1(n20856), .ip2(n20902), .ip3(n16776), .op(n16599) );
  and2_1 U18279 ( .ip1(n20735), .ip2(n16599), .op(n18748) );
  nand2_1 U18280 ( .ip1(n18927), .ip2(n20856), .op(n20894) );
  inv_1 U18281 ( .ip(n20894), .op(n20912) );
  inv_1 U18282 ( .ip(n19186), .op(n17523) );
  and2_1 U18283 ( .ip1(n16776), .ip2(n17575), .op(n20896) );
  nand3_1 U18284 ( .ip1(n20912), .ip2(n17523), .ip3(n20896), .op(n16600) );
  nand3_1 U18285 ( .ip1(n16601), .ip2(n18748), .ip3(n16600), .op(n16602) );
  ab_or_c_or_d U18286 ( .ip1(n16894), .ip2(n18374), .ip3(n16603), .ip4(n16602), 
        .op(n16604) );
  not_ab_or_c_or_d U18287 ( .ip1(n17529), .ip2(n20884), .ip3(n16605), .ip4(
        n16604), .op(n16615) );
  nand2_1 U18288 ( .ip1(n20892), .ip2(n12932), .op(n17489) );
  nand2_1 U18289 ( .ip1(n21536), .ip2(n10187), .op(n16607) );
  nand2_1 U18290 ( .ip1(n19056), .ip2(n10185), .op(n16606) );
  nand2_1 U18291 ( .ip1(n18927), .ip2(n13022), .op(n16766) );
  and4_1 U18292 ( .ip1(n17489), .ip2(n16607), .ip3(n16606), .ip4(n16766), .op(
        n16897) );
  mux2_1 U18293 ( .ip1(n13870), .ip2(n16608), .s(n21553), .op(n17478) );
  nor2_1 U18294 ( .ip1(n10184), .ip2(n17269), .op(n16609) );
  nor2_1 U18295 ( .ip1(n17492), .ip2(n21532), .op(n16758) );
  ab_or_c_or_d U18296 ( .ip1(n17478), .ip2(n16732), .ip3(n16609), .ip4(n16758), 
        .op(n16892) );
  mux2_1 U18297 ( .ip1(n16897), .ip2(n16892), .s(n10198), .op(n19423) );
  inv_1 U18298 ( .ip(n19423), .op(n17014) );
  nand2_1 U18299 ( .ip1(n17014), .ip2(n17547), .op(n16614) );
  nand2_1 U18300 ( .ip1(n20892), .ip2(n19068), .op(n18930) );
  nand2_1 U18301 ( .ip1(n18927), .ip2(n19199), .op(n19189) );
  mux2_1 U18302 ( .ip1(n20891), .ip2(n17073), .s(n21552), .op(n18914) );
  nand2_1 U18303 ( .ip1(n18914), .ip2(n17480), .op(n16611) );
  nand2_1 U18304 ( .ip1(n16610), .ip2(n16611), .op(n19204) );
  nand2_1 U18305 ( .ip1(n21536), .ip2(n16914), .op(n19190) );
  nand2_1 U18306 ( .ip1(n20892), .ip2(n10186), .op(n18364) );
  nand2_1 U18307 ( .ip1(n19056), .ip2(n19051), .op(n18929) );
  mux2_1 U18308 ( .ip1(n19204), .ip2(n16777), .s(n17575), .op(n19428) );
  nand2_1 U18309 ( .ip1(n19428), .ip2(n20736), .op(n16613) );
  nand2_1 U18310 ( .ip1(n16617), .ip2(n16827), .op(n16624) );
  inv_1 U18311 ( .ip(n16619), .op(n17255) );
  nor2_1 U18312 ( .ip1(n19419), .ip2(n17255), .op(n16618) );
  nor2_1 U18313 ( .ip1(n16880), .ip2(n16618), .op(n16622) );
  nand2_1 U18314 ( .ip1(n19417), .ip2(n16619), .op(n16620) );
  or2_1 U18315 ( .ip1(n16620), .ip2(n20717), .op(n16621) );
  nand2_1 U18316 ( .ip1(n16622), .ip2(n16621), .op(n16623) );
  xnor2_1 U18317 ( .ip1(n16624), .ip2(n16623), .op(n16625) );
  nand2_1 U18318 ( .ip1(n16625), .ip2(n21577), .op(n16664) );
  nand2_1 U18319 ( .ip1(n20892), .ip2(n16626), .op(n16685) );
  nand2_1 U18320 ( .ip1(n21536), .ip2(n19433), .op(n16629) );
  nand2_1 U18321 ( .ip1(n19056), .ip2(n12138), .op(n16628) );
  nand2_1 U18322 ( .ip1(n18927), .ip2(n16627), .op(n16658) );
  nand2_1 U18323 ( .ip1(n21536), .ip2(n10193), .op(n16631) );
  nand2_1 U18324 ( .ip1(n20892), .ip2(n16811), .op(n16630) );
  nand2_1 U18325 ( .ip1(n10206), .ip2(n18927), .op(n17450) );
  or2_1 U18326 ( .ip1(n12932), .ip2(n17267), .op(n16761) );
  nor2_1 U18327 ( .ip1(n18948), .ip2(n16873), .op(n16648) );
  inv_1 U18328 ( .ip(n17547), .op(n16893) );
  nor3_1 U18329 ( .ip1(n17443), .ip2(n16893), .ip3(n17478), .op(n16636) );
  nand2_1 U18330 ( .ip1(n16526), .ip2(n16632), .op(n16634) );
  nor3_1 U18331 ( .ip1(n16632), .ip2(n21551), .ip3(n16526), .op(n16633) );
  ab_or_c_or_d U18332 ( .ip1(n21557), .ip2(n16634), .ip3(n19066), .ip4(n16633), 
        .op(n16635) );
  not_ab_or_c_or_d U18333 ( .ip1(n20911), .ip2(n16637), .ip3(n16636), .ip4(
        n16635), .op(n16646) );
  nand2_1 U18334 ( .ip1(n21536), .ip2(n16423), .op(n16640) );
  nand2_1 U18335 ( .ip1(n18927), .ip2(n20221), .op(n16639) );
  nand2_1 U18336 ( .ip1(n20892), .ip2(n16838), .op(n16638) );
  nand2_1 U18337 ( .ip1(n19056), .ip2(n16973), .op(n16765) );
  nand2_1 U18338 ( .ip1(n18944), .ip2(n17529), .op(n16645) );
  nand2_1 U18339 ( .ip1(n21536), .ip2(n17492), .op(n16643) );
  nand2_1 U18340 ( .ip1(n18927), .ip2(n10187), .op(n17488) );
  nand2_1 U18341 ( .ip1(n20892), .ip2(n10185), .op(n16642) );
  nand2_1 U18342 ( .ip1(n19056), .ip2(n10184), .op(n16641) );
  nand2_1 U18343 ( .ip1(n17542), .ip2(n18374), .op(n16644) );
  nand3_1 U18344 ( .ip1(n16646), .ip2(n16645), .ip3(n16644), .op(n16647) );
  not_ab_or_c_or_d U18345 ( .ip1(n17541), .ip2(n18934), .ip3(n16648), .ip4(
        n16647), .op(n16663) );
  nor2_1 U18346 ( .ip1(n17267), .ip2(n10180), .op(n20890) );
  inv_1 U18347 ( .ip(n20890), .op(n16649) );
  nand2_1 U18348 ( .ip1(n20892), .ip2(n19051), .op(n19188) );
  nand2_1 U18349 ( .ip1(n18927), .ip2(n16914), .op(n18363) );
  nand2_1 U18350 ( .ip1(n21536), .ip2(n19199), .op(n18932) );
  nand2_1 U18351 ( .ip1(n17519), .ip2(n17575), .op(n16652) );
  inv_1 U18352 ( .ip(n17237), .op(n17034) );
  nand2_1 U18353 ( .ip1(n17034), .ip2(n20856), .op(n16651) );
  nand2_1 U18354 ( .ip1(n18914), .ip2(n17543), .op(n16650) );
  nand3_1 U18355 ( .ip1(n16652), .ip2(n16651), .ip3(n16650), .op(n17439) );
  inv_1 U18356 ( .ip(n17558), .op(n19205) );
  nand2_1 U18357 ( .ip1(n17439), .ip2(n19205), .op(n16656) );
  nand2_1 U18358 ( .ip1(n18914), .ip2(n17097), .op(n16654) );
  nand2_1 U18359 ( .ip1(n21536), .ip2(n20856), .op(n16653) );
  nand2_1 U18360 ( .ip1(n16654), .ip2(n16653), .op(n20229) );
  mux2_1 U18361 ( .ip1(n20229), .ip2(n17519), .s(n17575), .op(n17440) );
  nand2_1 U18362 ( .ip1(n17440), .ip2(n17523), .op(n16655) );
  nand2_1 U18363 ( .ip1(n16656), .ip2(n16655), .op(n18382) );
  nand2_1 U18364 ( .ip1(n18382), .ip2(n16776), .op(n16662) );
  nand2_1 U18365 ( .ip1(n19056), .ip2(n10186), .op(n19187) );
  nand2_1 U18366 ( .ip1(n21536), .ip2(n18738), .op(n18362) );
  nand2_1 U18367 ( .ip1(n18927), .ip2(n17530), .op(n17526) );
  nand2_1 U18368 ( .ip1(n21536), .ip2(n10188), .op(n17525) );
  mux2_1 U18369 ( .ip1(n17520), .ip2(n20230), .s(n17575), .op(n17467) );
  nand2_1 U18370 ( .ip1(n17467), .ip2(n20736), .op(n16661) );
  nand2_1 U18371 ( .ip1(n20715), .ip2(n20710), .op(n16668) );
  inv_1 U18372 ( .ip(n16665), .op(n20716) );
  nand2_1 U18373 ( .ip1(n20210), .ip2(n20716), .op(n16666) );
  nand2_1 U18374 ( .ip1(n20712), .ip2(n16666), .op(n16667) );
  xnor2_1 U18375 ( .ip1(n16668), .ip2(n16667), .op(n16669) );
  nand2_1 U18376 ( .ip1(n16669), .ip2(n21577), .op(n16703) );
  inv_1 U18377 ( .ip(n20239), .op(n17573) );
  inv_1 U18378 ( .ip(n19204), .op(n16674) );
  nor2_1 U18379 ( .ip1(n17573), .ip2(n16674), .op(n16671) );
  mux2_1 U18380 ( .ip1(n19066), .ip2(n16671), .s(n19427), .op(n16677) );
  inv_1 U18381 ( .ip(n16672), .op(n16673) );
  and2_1 U18382 ( .ip1(n17199), .ip2(n16673), .op(n19429) );
  inv_1 U18383 ( .ip(n19429), .op(n16675) );
  mux2_1 U18384 ( .ip1(n20894), .ip2(n16674), .s(n17575), .op(n19184) );
  nor3_1 U18385 ( .ip1(n16776), .ip2(n16675), .ip3(n19184), .op(n16676) );
  nor2_1 U18386 ( .ip1(n16677), .ip2(n16676), .op(n16702) );
  nand2_1 U18387 ( .ip1(n20892), .ip2(n17270), .op(n17527) );
  nand2_1 U18388 ( .ip1(n19056), .ip2(n18737), .op(n18361) );
  mux2_1 U18389 ( .ip1(n16777), .ip2(n19441), .s(n17575), .op(n16697) );
  nand2_1 U18390 ( .ip1(n21536), .ip2(n13678), .op(n16683) );
  nand2_1 U18391 ( .ip1(n13552), .ip2(n18927), .op(n16682) );
  nand2_1 U18392 ( .ip1(n20892), .ip2(n10189), .op(n16681) );
  nand2_1 U18393 ( .ip1(n16506), .ip2(n19056), .op(n16680) );
  nor2_1 U18394 ( .ip1(n10198), .ip2(n17498), .op(n19440) );
  inv_1 U18395 ( .ip(n19440), .op(n20218) );
  nor2_1 U18396 ( .ip1(n17001), .ip2(n20218), .op(n16696) );
  nor2_1 U18397 ( .ip1(n17575), .ip2(n17498), .op(n20231) );
  nand2_1 U18398 ( .ip1(n19056), .ip2(n16684), .op(n17524) );
  nand2_1 U18399 ( .ip1(n20231), .ip2(n19439), .op(n16694) );
  nand2_1 U18400 ( .ip1(n16688), .ip2(n20911), .op(n16693) );
  nand2_1 U18401 ( .ip1(n13552), .ip2(n13676), .op(n16689) );
  nand2_1 U18402 ( .ip1(n16689), .ip2(n21557), .op(n16692) );
  inv_1 U18403 ( .ip(n21551), .op(n20904) );
  nand3_1 U18404 ( .ip1(n16423), .ip2(n20904), .ip3(n16690), .op(n16691) );
  not_ab_or_c_or_d U18405 ( .ip1(n21549), .ip2(n16697), .ip3(n16696), .ip4(
        n16695), .op(n16701) );
  inv_1 U18406 ( .ip(n20896), .op(n18936) );
  nor2_1 U18407 ( .ip1(n18936), .ip2(n16892), .op(n16699) );
  nor2_1 U18408 ( .ip1(n17575), .ip2(n16776), .op(n21540) );
  inv_1 U18409 ( .ip(n21540), .op(n20887) );
  nor2_1 U18410 ( .ip1(n20887), .ip2(n16897), .op(n16698) );
  ab_or_c_or_d U18411 ( .ip1(n16894), .ip2(n19427), .ip3(n16699), .ip4(n16698), 
        .op(n19212) );
  inv_1 U18412 ( .ip(n20724), .op(n20900) );
  nand2_1 U18413 ( .ip1(n19212), .ip2(n20900), .op(n16700) );
  inv_1 U18414 ( .ip(n16704), .op(n17505) );
  nand2_1 U18415 ( .ip1(n17503), .ip2(n17505), .op(n16705) );
  nand2_1 U18416 ( .ip1(n17504), .ip2(n16705), .op(n16710) );
  inv_1 U18417 ( .ip(n16706), .op(n16708) );
  nand2_1 U18418 ( .ip1(n16708), .ip2(n16707), .op(n16709) );
  xnor2_1 U18419 ( .ip1(n16710), .ip2(n16709), .op(n16711) );
  nand2_1 U18420 ( .ip1(n16711), .ip2(n21577), .op(n16749) );
  inv_1 U18421 ( .ip(n17443), .op(n18913) );
  nand2_1 U18422 ( .ip1(n17035), .ip2(n18913), .op(n16713) );
  inv_1 U18423 ( .ip(n21534), .op(n17236) );
  inv_1 U18424 ( .ip(n17223), .op(n17493) );
  nand2_1 U18425 ( .ip1(n17236), .ip2(n17493), .op(n16712) );
  nand2_1 U18426 ( .ip1(n16713), .ip2(n16712), .op(n16954) );
  nor2_1 U18427 ( .ip1(n10198), .ip2(n10184), .op(n16714) );
  nor2_1 U18428 ( .ip1(n20907), .ip2(n16714), .op(n16716) );
  nor3_1 U18429 ( .ip1(n17575), .ip2(n21551), .ip3(n13728), .op(n16715) );
  ab_or_c_or_d U18430 ( .ip1(n16717), .ip2(n20911), .ip3(n16716), .ip4(n16715), 
        .op(n16723) );
  or2_1 U18431 ( .ip1(n20239), .ip2(n19429), .op(n21544) );
  nand2_1 U18432 ( .ip1(n21544), .ip2(n13881), .op(n21565) );
  nor2_1 U18433 ( .ip1(n17237), .ip2(n17226), .op(n16721) );
  nor2_1 U18434 ( .ip1(n17443), .ip2(n17208), .op(n16720) );
  nor2_1 U18435 ( .ip1(n17223), .ip2(n17225), .op(n16719) );
  nor2_1 U18436 ( .ip1(n17227), .ip2(n17222), .op(n16718) );
  or4_1 U18437 ( .ip1(n16721), .ip2(n16720), .ip3(n16719), .ip4(n16718), .op(
        n16969) );
  nor2_1 U18438 ( .ip1(n21565), .ip2(n16969), .op(n16722) );
  not_ab_or_c_or_d U18439 ( .ip1(n21562), .ip2(n16954), .ip3(n16723), .ip4(
        n16722), .op(n16748) );
  nand2_1 U18440 ( .ip1(n21536), .ip2(n10180), .op(n16725) );
  nand2_1 U18441 ( .ip1(n10191), .ip2(n19056), .op(n16724) );
  nand2_1 U18442 ( .ip1(n16725), .ip2(n16724), .op(n16727) );
  nor2_1 U18443 ( .ip1(n13525), .ip2(n17224), .op(n16726) );
  nor2_1 U18444 ( .ip1(n16727), .ip2(n16726), .op(n17058) );
  nand2_1 U18445 ( .ip1(n17058), .ip2(n17575), .op(n16729) );
  nand2_1 U18446 ( .ip1(n17121), .ip2(n17543), .op(n16728) );
  nand2_1 U18447 ( .ip1(n16729), .ip2(n16728), .op(n16957) );
  nand2_1 U18448 ( .ip1(n16957), .ip2(n21544), .op(n16731) );
  inv_1 U18449 ( .ip(n20856), .op(n20905) );
  nor3_1 U18450 ( .ip1(n17097), .ip2(n17575), .ip3(n20905), .op(n16859) );
  nand2_1 U18451 ( .ip1(n16859), .ip2(n20239), .op(n16730) );
  nand2_1 U18452 ( .ip1(n16731), .ip2(n16730), .op(n16981) );
  nand2_1 U18453 ( .ip1(n16981), .ip2(n16776), .op(n16747) );
  mux2_1 U18454 ( .ip1(n13678), .ip2(n10189), .s(n21553), .op(n16806) );
  nand2_1 U18455 ( .ip1(n16806), .ip2(n16732), .op(n16734) );
  nand2_1 U18456 ( .ip1(n13877), .ip2(n18927), .op(n16868) );
  nand3_1 U18457 ( .ip1(n16734), .ip2(n16733), .ip3(n16868), .op(n17055) );
  nor2_1 U18458 ( .ip1(n17237), .ip2(n17207), .op(n16736) );
  mux2_1 U18459 ( .ip1(n12138), .ip2(n19433), .s(n21552), .op(n17209) );
  nor2_1 U18460 ( .ip1(n17227), .ip2(n17209), .op(n16735) );
  not_ab_or_c_or_d U18461 ( .ip1(n17575), .ip2(n17055), .ip3(n16736), .ip4(
        n16735), .op(n16980) );
  or2_1 U18462 ( .ip1(n13166), .ip2(n16980), .op(n16745) );
  nand2_1 U18463 ( .ip1(n21536), .ip2(n16811), .op(n16869) );
  nand2_1 U18464 ( .ip1(n17042), .ip2(n18927), .op(n16851) );
  nand4_1 U18465 ( .ip1(n16738), .ip2(n16737), .ip3(n16869), .ip4(n16851), 
        .op(n17047) );
  nand2_1 U18466 ( .ip1(n17047), .ip2(n21540), .op(n16744) );
  nor2_1 U18467 ( .ip1(n10195), .ip2(n17269), .op(n16739) );
  not_ab_or_c_or_d U18468 ( .ip1(n21536), .ip2(n10185), .ip3(n18918), .ip4(
        n16739), .op(n16742) );
  nand2_1 U18469 ( .ip1(n18927), .ip2(n10184), .op(n16741) );
  nand2_1 U18470 ( .ip1(n19056), .ip2(n10187), .op(n16740) );
  nand3_1 U18471 ( .ip1(n16742), .ip2(n16741), .ip3(n16740), .op(n16743) );
  nand4_1 U18472 ( .ip1(n16745), .ip2(n21572), .ip3(n16744), .ip4(n16743), 
        .op(n16746) );
  inv_1 U18473 ( .ip(n17193), .op(n16751) );
  nand2_1 U18474 ( .ip1(n16751), .ip2(n16750), .op(n16752) );
  inv_1 U18475 ( .ip(n17565), .op(n17024) );
  xnor2_1 U18476 ( .ip1(n16752), .ip2(n17024), .op(n16753) );
  nand2_1 U18477 ( .ip1(n16753), .ip2(n21577), .op(n16787) );
  inv_1 U18478 ( .ip(n16892), .op(n16775) );
  nand2_1 U18479 ( .ip1(n10195), .ip2(n13881), .op(n16757) );
  nor3_1 U18480 ( .ip1(n13166), .ip2(n21551), .ip3(n10195), .op(n16756) );
  nor2_1 U18481 ( .ip1(n21555), .ip2(n16754), .op(n16755) );
  ab_or_c_or_d U18482 ( .ip1(n21557), .ip2(n16757), .ip3(n16756), .ip4(n16755), 
        .op(n16774) );
  inv_1 U18483 ( .ip(n16758), .op(n16762) );
  nand2_1 U18484 ( .ip1(n21536), .ip2(n16446), .op(n16760) );
  nand2_1 U18485 ( .ip1(n20892), .ip2(n13540), .op(n16759) );
  inv_1 U18486 ( .ip(n19193), .op(n20885) );
  nor2_1 U18487 ( .ip1(n20885), .ip2(n19439), .op(n16771) );
  inv_1 U18488 ( .ip(n16763), .op(n16767) );
  nand2_1 U18489 ( .ip1(n20892), .ip2(n13698), .op(n16764) );
  and4_1 U18490 ( .ip1(n16767), .ip2(n16766), .ip3(n16765), .ip4(n16764), .op(
        n16999) );
  nand2_1 U18491 ( .ip1(n16999), .ip2(n21540), .op(n16769) );
  nand2_1 U18492 ( .ip1(n17001), .ip2(n20896), .op(n16768) );
  nand3_1 U18493 ( .ip1(n16769), .ip2(n21572), .ip3(n16768), .op(n16770) );
  not_ab_or_c_or_d U18494 ( .ip1(n19427), .ip2(n16772), .ip3(n16771), .ip4(
        n16770), .op(n16773) );
  not_ab_or_c_or_d U18495 ( .ip1(n17541), .ip2(n16775), .ip3(n16774), .ip4(
        n16773), .op(n16786) );
  nand2_1 U18496 ( .ip1(n19184), .ip2(n16776), .op(n16780) );
  nor2_1 U18497 ( .ip1(n20887), .ip2(n16777), .op(n16779) );
  nor2_1 U18498 ( .ip1(n18918), .ip2(n19441), .op(n16778) );
  nor2_1 U18499 ( .ip1(n16779), .ip2(n16778), .op(n16781) );
  and2_1 U18500 ( .ip1(n16780), .ip2(n16781), .op(n16906) );
  nand2_1 U18501 ( .ip1(n16906), .ip2(n19429), .op(n16785) );
  nor2_1 U18502 ( .ip1(n18936), .ip2(n19204), .op(n16783) );
  inv_1 U18503 ( .ip(n16781), .op(n16782) );
  not_ab_or_c_or_d U18504 ( .ip1(n20905), .ip2(n19193), .ip3(n16783), .ip4(
        n16782), .op(n16907) );
  nand2_1 U18505 ( .ip1(n16907), .ip2(n20239), .op(n16784) );
  inv_1 U18506 ( .ip(n16987), .op(n16793) );
  nor2_1 U18507 ( .ip1(n16995), .ip2(n16791), .op(n16792) );
  nor2_1 U18508 ( .ip1(n16793), .ip2(n16792), .op(n16799) );
  nand2_1 U18509 ( .ip1(n16990), .ip2(n16988), .op(n16795) );
  inv_1 U18510 ( .ip(n17567), .op(n17026) );
  or2_1 U18511 ( .ip1(n16795), .ip2(n17026), .op(n16798) );
  inv_1 U18512 ( .ip(n16794), .op(n17564) );
  nor2_1 U18513 ( .ip1(n17564), .ip2(n16795), .op(n16796) );
  nand2_1 U18514 ( .ip1(n16796), .ip2(n17024), .op(n16797) );
  nand3_1 U18515 ( .ip1(n16799), .ip2(n16798), .ip3(n16797), .op(n16800) );
  xnor2_1 U18516 ( .ip1(n16790), .ip2(n16800), .op(n16801) );
  inv_1 U18517 ( .ip(n16801), .op(n16802) );
  nand2_1 U18518 ( .ip1(n16802), .ip2(n21577), .op(n16823) );
  nand2_1 U18519 ( .ip1(n20892), .ip2(n10206), .op(n16867) );
  nand2_1 U18520 ( .ip1(n13552), .ip2(n19056), .op(n16803) );
  nand4_1 U18521 ( .ip1(n16805), .ip2(n16804), .ip3(n16867), .ip4(n16803), 
        .op(n17201) );
  nor2_1 U18522 ( .ip1(n17237), .ip2(n17209), .op(n16808) );
  inv_1 U18523 ( .ip(n16806), .op(n17210) );
  nor2_1 U18524 ( .ip1(n17227), .ip2(n17210), .op(n16807) );
  not_ab_or_c_or_d U18525 ( .ip1(n17575), .ip2(n17201), .ip3(n16808), .ip4(
        n16807), .op(n21550) );
  inv_1 U18526 ( .ip(n21549), .op(n20726) );
  nor2_1 U18527 ( .ip1(n20726), .ip2(n21564), .op(n16817) );
  or2_1 U18528 ( .ip1(n13166), .ip2(n20735), .op(n17462) );
  inv_1 U18529 ( .ip(n16809), .op(n16810) );
  nand2_1 U18530 ( .ip1(n16810), .ip2(n20911), .op(n16815) );
  nand2_1 U18531 ( .ip1(n16811), .ip2(n13702), .op(n16812) );
  nand2_1 U18532 ( .ip1(n16812), .ip2(n21557), .op(n16814) );
  nand3_1 U18533 ( .ip1(n13698), .ip2(n20904), .ip3(n12596), .op(n16813) );
  not_ab_or_c_or_d U18534 ( .ip1(n20736), .ip2(n21550), .ip3(n16817), .ip4(
        n16816), .op(n16822) );
  nand2_1 U18535 ( .ip1(n18913), .ip2(n16776), .op(n17554) );
  nor2_1 U18536 ( .ip1(n21534), .ip2(n17554), .op(n16819) );
  nor2_1 U18537 ( .ip1(n18918), .ip2(n19050), .op(n16818) );
  not_ab_or_c_or_d U18538 ( .ip1(n21540), .ip2(n17235), .ip3(n16819), .ip4(
        n16818), .op(n18728) );
  or2_1 U18539 ( .ip1(n20724), .ip2(n18728), .op(n16821) );
  inv_1 U18540 ( .ip(n21565), .op(n17015) );
  nand2_1 U18541 ( .ip1(n18729), .ip2(n17015), .op(n16820) );
  nand2_1 U18542 ( .ip1(n16825), .ip2(n16824), .op(n16836) );
  inv_1 U18543 ( .ip(n16880), .op(n17252) );
  or2_1 U18544 ( .ip1(n16828), .ip2(n17252), .op(n16826) );
  nand2_1 U18545 ( .ip1(n16827), .ip2(n16826), .op(n16830) );
  nor2_1 U18546 ( .ip1(n17255), .ip2(n16828), .op(n16831) );
  inv_1 U18547 ( .ip(n19419), .op(n17257) );
  and2_1 U18548 ( .ip1(n16831), .ip2(n17257), .op(n16829) );
  nor2_1 U18549 ( .ip1(n16830), .ip2(n16829), .op(n16834) );
  nand2_1 U18550 ( .ip1(n19417), .ip2(n16831), .op(n16832) );
  or2_1 U18551 ( .ip1(n16832), .ip2(n20717), .op(n16833) );
  nand2_1 U18552 ( .ip1(n16834), .ip2(n16833), .op(n16835) );
  xnor2_1 U18553 ( .ip1(n16836), .ip2(n16835), .op(n16837) );
  nand2_1 U18554 ( .ip1(n16837), .ip2(n21577), .op(n16879) );
  nand2_1 U18555 ( .ip1(n21536), .ip2(n16838), .op(n16840) );
  nand2_1 U18556 ( .ip1(n18927), .ip2(n12138), .op(n16839) );
  nand2_1 U18557 ( .ip1(n16840), .ip2(n16839), .op(n16844) );
  nand2_1 U18558 ( .ip1(n20892), .ip2(n20221), .op(n16842) );
  nand2_1 U18559 ( .ip1(n19056), .ip2(n16423), .op(n16841) );
  nand2_1 U18560 ( .ip1(n16842), .ip2(n16841), .op(n16843) );
  nor2_1 U18561 ( .ip1(n16844), .ip2(n16843), .op(n17120) );
  inv_1 U18562 ( .ip(n17120), .op(n17170) );
  nand2_1 U18563 ( .ip1(n21536), .ip2(n16845), .op(n16850) );
  nand2_1 U18564 ( .ip1(n18927), .ip2(n16854), .op(n16849) );
  nand2_1 U18565 ( .ip1(n20892), .ip2(n16627), .op(n16848) );
  nand2_1 U18566 ( .ip1(n19056), .ip2(n16846), .op(n16847) );
  inv_1 U18567 ( .ip(n17166), .op(n17115) );
  nor2_1 U18568 ( .ip1(n17275), .ip2(n17115), .op(n16865) );
  nand2_1 U18569 ( .ip1(n20892), .ip2(n16446), .op(n16853) );
  nand2_1 U18570 ( .ip1(n21536), .ip2(n13540), .op(n16852) );
  or2_1 U18571 ( .ip1(n17492), .ip2(n17267), .op(n21537) );
  inv_1 U18572 ( .ip(n18374), .op(n17528) );
  or2_1 U18573 ( .ip1(n17033), .ip2(n17528), .op(n16863) );
  nand2_1 U18574 ( .ip1(n10190), .ip2(n16855), .op(n16857) );
  nor3_1 U18575 ( .ip1(n16855), .ip2(n21551), .ip3(n10190), .op(n16856) );
  not_ab_or_c_or_d U18576 ( .ip1(n21557), .ip2(n16857), .ip3(n16856), .ip4(
        n19066), .op(n16862) );
  nand2_1 U18577 ( .ip1(n16858), .ip2(n20911), .op(n16861) );
  nand2_1 U18578 ( .ip1(n16859), .ip2(n19205), .op(n16931) );
  or2_1 U18579 ( .ip1(n13166), .ip2(n16931), .op(n16860) );
  not_ab_or_c_or_d U18580 ( .ip1(n17529), .ip2(n17170), .ip3(n16865), .ip4(
        n16864), .op(n16878) );
  nand2_1 U18581 ( .ip1(n10193), .ip2(n19056), .op(n16866) );
  nand2_1 U18582 ( .ip1(n16867), .ip2(n16866), .op(n16871) );
  nand2_1 U18583 ( .ip1(n16869), .ip2(n16868), .op(n16870) );
  nor2_1 U18584 ( .ip1(n16871), .ip2(n16870), .op(n17178) );
  inv_1 U18585 ( .ip(n17178), .op(n16872) );
  nor2_1 U18586 ( .ip1(n16873), .ip2(n16872), .op(n16875) );
  nor2_1 U18587 ( .ip1(n17498), .ip2(n16969), .op(n16874) );
  not_ab_or_c_or_d U18588 ( .ip1(n17547), .ip2(n16954), .ip3(n16875), .ip4(
        n16874), .op(n16877) );
  nand2_1 U18589 ( .ip1(n16957), .ip2(n21549), .op(n16876) );
  nand2_1 U18590 ( .ip1(n17250), .ip2(n17245), .op(n16890) );
  inv_1 U18591 ( .ip(n16882), .op(n17251) );
  nand2_1 U18592 ( .ip1(n16880), .ip2(n17251), .op(n16881) );
  nand2_1 U18593 ( .ip1(n17247), .ip2(n16881), .op(n16884) );
  nor2_1 U18594 ( .ip1(n17255), .ip2(n16882), .op(n16885) );
  and2_1 U18595 ( .ip1(n16885), .ip2(n17257), .op(n16883) );
  nor2_1 U18596 ( .ip1(n16884), .ip2(n16883), .op(n16888) );
  nand2_1 U18597 ( .ip1(n19417), .ip2(n16885), .op(n16886) );
  or2_1 U18598 ( .ip1(n16886), .ip2(n20717), .op(n16887) );
  nand2_1 U18599 ( .ip1(n16888), .ip2(n16887), .op(n16889) );
  xnor2_1 U18600 ( .ip1(n16890), .ip2(n16889), .op(n16891) );
  nand2_1 U18601 ( .ip1(n16891), .ip2(n21577), .op(n16911) );
  nor3_1 U18602 ( .ip1(n10198), .ip2(n16893), .ip3(n16892), .op(n16905) );
  nand2_1 U18603 ( .ip1(n16894), .ip2(n18367), .op(n16903) );
  nand2_1 U18604 ( .ip1(n10517), .ip2(n10197), .op(n16896) );
  nor3_1 U18605 ( .ip1(n10197), .ip2(n21551), .ip3(n10517), .op(n16895) );
  ab_or_c_or_d U18606 ( .ip1(n21557), .ip2(n16896), .ip3(n19066), .ip4(n16895), 
        .op(n16899) );
  nor2_1 U18607 ( .ip1(n17528), .ip2(n16897), .op(n16898) );
  not_ab_or_c_or_d U18608 ( .ip1(n20911), .ip2(n16900), .ip3(n16899), .ip4(
        n16898), .op(n16902) );
  nand2_1 U18609 ( .ip1(n20884), .ip2(n17541), .op(n16901) );
  nand3_1 U18610 ( .ip1(n16903), .ip2(n16902), .ip3(n16901), .op(n16904) );
  not_ab_or_c_or_d U18611 ( .ip1(n17529), .ip2(n19426), .ip3(n16905), .ip4(
        n16904), .op(n16910) );
  nand2_1 U18612 ( .ip1(n16906), .ip2(n17523), .op(n16909) );
  nand2_1 U18613 ( .ip1(n16907), .ip2(n19205), .op(n16908) );
  xor2_1 U18614 ( .ip1(n16935), .ip2(n20855), .op(n16912) );
  nor2_1 U18615 ( .ip1(n16912), .ip2(n19051), .op(n19172) );
  inv_1 U18616 ( .ip(n19172), .op(n19175) );
  nand2_1 U18617 ( .ip1(n16912), .ip2(n19051), .op(n17081) );
  nand2_1 U18618 ( .ip1(n19175), .ip2(n17081), .op(n16929) );
  xor2_1 U18619 ( .ip1(n18369), .ip2(n16913), .op(n16915) );
  nand2_1 U18620 ( .ip1(n16915), .ip2(n16914), .op(n18349) );
  nor2_1 U18621 ( .ip1(n16915), .ip2(n16914), .op(n16921) );
  inv_1 U18622 ( .ip(n16921), .op(n18350) );
  xor2_1 U18623 ( .ip1(n18731), .ip2(n20855), .op(n16920) );
  nand2_1 U18624 ( .ip1(n16920), .ip2(n10186), .op(n18721) );
  inv_1 U18625 ( .ip(n18721), .op(n18353) );
  nand2_1 U18626 ( .ip1(n18350), .ip2(n18353), .op(n16916) );
  nand2_1 U18627 ( .ip1(n18349), .ip2(n16916), .op(n16923) );
  or2_1 U18628 ( .ip1(n16924), .ip2(n16917), .op(n16918) );
  nand2_1 U18629 ( .ip1(n16919), .ip2(n16918), .op(n18351) );
  nor2_1 U18630 ( .ip1(n16920), .ip2(n10186), .op(n18354) );
  nor2_1 U18631 ( .ip1(n18354), .ip2(n16921), .op(n16926) );
  and2_1 U18632 ( .ip1(n18351), .ip2(n16926), .op(n16922) );
  nor2_1 U18633 ( .ip1(n16923), .ip2(n16922), .op(n20871) );
  nor2_1 U18634 ( .ip1(n16925), .ip2(n16924), .op(n18723) );
  nand2_1 U18635 ( .ip1(n18723), .ip2(n16926), .op(n20876) );
  inv_1 U18636 ( .ip(n20876), .op(n19176) );
  nand2_1 U18637 ( .ip1(n20878), .ip2(n19176), .op(n16927) );
  nand2_1 U18638 ( .ip1(n20871), .ip2(n16927), .op(n16928) );
  xnor2_1 U18639 ( .ip1(n16929), .ip2(n16928), .op(n16930) );
  nand2_1 U18640 ( .ip1(n16930), .ip2(n21577), .op(n16961) );
  nand2_1 U18641 ( .ip1(n19205), .ip2(n20856), .op(n19064) );
  inv_1 U18642 ( .ip(n19064), .op(n16953) );
  nand2_1 U18643 ( .ip1(n16931), .ip2(n13166), .op(n16952) );
  nand2_1 U18644 ( .ip1(n16932), .ip2(n20911), .op(n16938) );
  nand2_1 U18645 ( .ip1(n10178), .ip2(n16933), .op(n16934) );
  nand2_1 U18646 ( .ip1(n16934), .ip2(n21557), .op(n16937) );
  nand3_1 U18647 ( .ip1(n19051), .ip2(n20904), .ip3(n16935), .op(n16936) );
  nand4_1 U18648 ( .ip1(n16938), .ip2(n20735), .ip3(n16937), .ip4(n16936), 
        .op(n16951) );
  nand2_1 U18649 ( .ip1(n21536), .ip2(n17270), .op(n16942) );
  nand2_1 U18650 ( .ip1(n18927), .ip2(n18737), .op(n16941) );
  nand2_1 U18651 ( .ip1(n20892), .ip2(n17530), .op(n16940) );
  nand2_1 U18652 ( .ip1(n19056), .ip2(n10188), .op(n16939) );
  nor2_1 U18653 ( .ip1(n20887), .ip2(n17167), .op(n16949) );
  nor2_1 U18654 ( .ip1(n10178), .ip2(n21532), .op(n16946) );
  nor2_1 U18655 ( .ip1(n17267), .ip2(n13654), .op(n16945) );
  nor2_1 U18656 ( .ip1(n13656), .ip2(n17268), .op(n16944) );
  nor2_1 U18657 ( .ip1(n11941), .ip2(n17269), .op(n16943) );
  nor2_1 U18658 ( .ip1(n18936), .ip2(n17166), .op(n16947) );
  ab_or_c_or_d U18659 ( .ip1(n17106), .ip2(n19427), .ip3(n16947), .ip4(n20724), 
        .op(n16948) );
  not_ab_or_c_or_d U18660 ( .ip1(n17120), .ip2(n19193), .ip3(n16949), .ip4(
        n16948), .op(n16950) );
  not_ab_or_c_or_d U18661 ( .ip1(n16953), .ip2(n16952), .ip3(n16951), .ip4(
        n16950), .op(n16960) );
  nor2_1 U18662 ( .ip1(n13166), .ip2(n16954), .op(n16956) );
  nor2_1 U18663 ( .ip1(n18918), .ip2(n17178), .op(n16955) );
  not_ab_or_c_or_d U18664 ( .ip1(n21540), .ip2(n17033), .ip3(n16956), .ip4(
        n16955), .op(n16982) );
  inv_1 U18665 ( .ip(n20883), .op(n19213) );
  nand2_1 U18666 ( .ip1(n16982), .ip2(n19213), .op(n16959) );
  nand2_1 U18667 ( .ip1(n16957), .ip2(n20736), .op(n16958) );
  nand2_1 U18668 ( .ip1(n16963), .ip2(n16962), .op(n16967) );
  or2_1 U18669 ( .ip1(n16964), .ip2(n20717), .op(n16965) );
  nand2_1 U18670 ( .ip1(n17468), .ip2(n16965), .op(n16966) );
  xnor2_1 U18671 ( .ip1(n16967), .ip2(n16966), .op(n16968) );
  nand2_1 U18672 ( .ip1(n16968), .ip2(n21577), .op(n16986) );
  nor2_1 U18673 ( .ip1(n20726), .ip2(n16969), .op(n16979) );
  inv_1 U18674 ( .ip(n16970), .op(n16971) );
  or2_1 U18675 ( .ip1(n16971), .ip2(n21555), .op(n16977) );
  nand3_1 U18676 ( .ip1(n16973), .ip2(n20904), .ip3(n16972), .op(n16976) );
  nand2_1 U18677 ( .ip1(n13553), .ip2(n13708), .op(n16974) );
  nand2_1 U18678 ( .ip1(n16974), .ip2(n21557), .op(n16975) );
  not_ab_or_c_or_d U18679 ( .ip1(n20736), .ip2(n16980), .ip3(n16979), .ip4(
        n16978), .op(n16985) );
  nand2_1 U18680 ( .ip1(n16981), .ip2(n13166), .op(n16984) );
  nand2_1 U18681 ( .ip1(n16982), .ip2(n20900), .op(n16983) );
  nand2_1 U18682 ( .ip1(n17567), .ip2(n16990), .op(n16994) );
  nor2_1 U18683 ( .ip1(n17564), .ip2(n16991), .op(n16992) );
  nand2_1 U18684 ( .ip1(n17024), .ip2(n16992), .op(n16993) );
  nand3_1 U18685 ( .ip1(n16995), .ip2(n16994), .ip3(n16993), .op(n16996) );
  xnor2_1 U18686 ( .ip1(n16989), .ip2(n16996), .op(n16997) );
  inv_1 U18687 ( .ip(n16997), .op(n16998) );
  nand2_1 U18688 ( .ip1(n16998), .ip2(n21577), .op(n17019) );
  nand2_1 U18689 ( .ip1(n16999), .ip2(n19427), .op(n17005) );
  inv_1 U18690 ( .ip(n21572), .op(n17583) );
  nor2_1 U18691 ( .ip1(n20885), .ip2(n19441), .op(n17000) );
  not_ab_or_c_or_d U18692 ( .ip1(n21540), .ip2(n17001), .ip3(n17583), .ip4(
        n17000), .op(n17004) );
  inv_1 U18693 ( .ip(n19439), .op(n17002) );
  nand2_1 U18694 ( .ip1(n17002), .ip2(n20896), .op(n17003) );
  nand3_1 U18695 ( .ip1(n17005), .ip2(n17004), .ip3(n17003), .op(n17013) );
  nor3_1 U18696 ( .ip1(n17006), .ip2(n21551), .ip3(n10193), .op(n17009) );
  nor2_1 U18697 ( .ip1(n20907), .ip2(n17007), .op(n17008) );
  not_ab_or_c_or_d U18698 ( .ip1(n20911), .ip2(n17010), .ip3(n17009), .ip4(
        n17008), .op(n17012) );
  nand3_1 U18699 ( .ip1(n20912), .ip2(n20896), .ip3(n19429), .op(n17011) );
  and4_1 U18700 ( .ip1(n17013), .ip2(n17012), .ip3(n17462), .ip4(n17011), .op(
        n17018) );
  nand2_1 U18701 ( .ip1(n17014), .ip2(n21562), .op(n17017) );
  nand2_1 U18702 ( .ip1(n19428), .ip2(n17015), .op(n17016) );
  inv_1 U18703 ( .ip(n17020), .op(n17022) );
  nor2_1 U18704 ( .ip1(n17564), .ip2(n17561), .op(n17025) );
  nand2_1 U18705 ( .ip1(n17025), .ip2(n17024), .op(n17029) );
  or2_1 U18706 ( .ip1(n17561), .ip2(n17026), .op(n17027) );
  nand2_1 U18707 ( .ip1(n17029), .ip2(n17028), .op(n17030) );
  xnor2_1 U18708 ( .ip1(n17023), .ip2(n17030), .op(n17031) );
  inv_1 U18709 ( .ip(n17031), .op(n17032) );
  nand2_1 U18710 ( .ip1(n21577), .ip2(n17032), .op(n17072) );
  nand2_1 U18711 ( .ip1(n17033), .ip2(n17575), .op(n17039) );
  and2_1 U18712 ( .ip1(n21534), .ip2(n17034), .op(n17037) );
  nor2_1 U18713 ( .ip1(n17227), .ip2(n17035), .op(n17036) );
  nor2_1 U18714 ( .ip1(n17037), .ip2(n17036), .op(n17038) );
  and2_1 U18715 ( .ip1(n17039), .ip2(n17038), .op(n17184) );
  nor2_1 U18716 ( .ip1(n17040), .ip2(n12932), .op(n17041) );
  nor2_1 U18717 ( .ip1(n20907), .ip2(n17041), .op(n17045) );
  nor3_1 U18718 ( .ip1(n17043), .ip2(n21551), .ip3(n17042), .op(n17044) );
  ab_or_c_or_d U18719 ( .ip1(n17046), .ip2(n20911), .ip3(n17045), .ip4(n17044), 
        .op(n17057) );
  nand2_1 U18720 ( .ip1(n17047), .ip2(n19427), .op(n17048) );
  nand2_1 U18721 ( .ip1(n17048), .ip2(n21572), .op(n17054) );
  nor2_1 U18722 ( .ip1(n17237), .ip2(n17225), .op(n17052) );
  nor2_1 U18723 ( .ip1(n17227), .ip2(n17208), .op(n17051) );
  nor2_1 U18724 ( .ip1(n17443), .ip2(n17209), .op(n17050) );
  nor2_1 U18725 ( .ip1(n17223), .ip2(n17207), .op(n17049) );
  nor2_1 U18726 ( .ip1(n20736), .ip2(n17152), .op(n17053) );
  not_ab_or_c_or_d U18727 ( .ip1(n21540), .ip2(n17055), .ip3(n17054), .ip4(
        n17053), .op(n17056) );
  not_ab_or_c_or_d U18728 ( .ip1(n21562), .ip2(n17184), .ip3(n17057), .ip4(
        n17056), .op(n17071) );
  nand2_1 U18729 ( .ip1(n17443), .ip2(n20856), .op(n18916) );
  or2_1 U18730 ( .ip1(n17575), .ip2(n17058), .op(n17062) );
  nor2_1 U18731 ( .ip1(n17223), .ip2(n17226), .op(n17060) );
  nor2_1 U18732 ( .ip1(n17443), .ip2(n17222), .op(n17059) );
  nor2_1 U18733 ( .ip1(n17060), .ip2(n17059), .op(n17061) );
  nand2_1 U18734 ( .ip1(n17062), .ip2(n17061), .op(n17149) );
  mux2_1 U18735 ( .ip1(n18916), .ip2(n17149), .s(n13881), .op(n17065) );
  inv_1 U18736 ( .ip(n17554), .op(n17063) );
  nand2_1 U18737 ( .ip1(n17121), .ip2(n17063), .op(n17064) );
  nand2_1 U18738 ( .ip1(n17065), .ip2(n17064), .op(n17185) );
  nand2_1 U18739 ( .ip1(n17185), .ip2(n20239), .op(n17070) );
  inv_1 U18740 ( .ip(n17149), .op(n17066) );
  nand2_1 U18741 ( .ip1(n17066), .ip2(n13881), .op(n17068) );
  nand3_1 U18742 ( .ip1(n17121), .ip2(n17097), .ip3(n20896), .op(n17067) );
  nand2_1 U18743 ( .ip1(n17068), .ip2(n17067), .op(n17186) );
  nand2_1 U18744 ( .ip1(n17186), .ip2(n19429), .op(n17069) );
  xor2_1 U18745 ( .ip1(n17102), .ip2(n20855), .op(n17074) );
  nor2_1 U18746 ( .ip1(n17074), .ip2(n17073), .op(n20864) );
  inv_1 U18747 ( .ip(n20864), .op(n20860) );
  nand2_1 U18748 ( .ip1(n17074), .ip2(n17073), .op(n20863) );
  nand2_1 U18749 ( .ip1(n20860), .ip2(n20863), .op(n17095) );
  xor2_1 U18750 ( .ip1(n18920), .ip2(n20855), .op(n17075) );
  nand2_1 U18751 ( .ip1(n17075), .ip2(n20891), .op(n18902) );
  inv_1 U18752 ( .ip(n18902), .op(n17077) );
  nor2_1 U18753 ( .ip1(n17075), .ip2(n20891), .op(n17079) );
  xor2_1 U18754 ( .ip1(n20855), .ip2(n19069), .op(n17078) );
  nand2_1 U18755 ( .ip1(n17078), .ip2(n19068), .op(n19040) );
  nor2_1 U18756 ( .ip1(n17079), .ip2(n19040), .op(n17076) );
  or2_1 U18757 ( .ip1(n17077), .ip2(n17076), .op(n20861) );
  nor2_1 U18758 ( .ip1(n17078), .ip2(n19068), .op(n18904) );
  inv_1 U18759 ( .ip(n18904), .op(n19041) );
  inv_1 U18760 ( .ip(n17079), .op(n18903) );
  nand2_1 U18761 ( .ip1(n19041), .ip2(n18903), .op(n20865) );
  xor2_1 U18762 ( .ip1(n13601), .ip2(n20855), .op(n17080) );
  nand2_1 U18763 ( .ip1(n17080), .ip2(n19199), .op(n19170) );
  nor2_1 U18764 ( .ip1(n17080), .ip2(n19199), .op(n17083) );
  inv_1 U18765 ( .ip(n17083), .op(n19171) );
  inv_1 U18766 ( .ip(n17081), .op(n19174) );
  nand2_1 U18767 ( .ip1(n19171), .ip2(n19174), .op(n17082) );
  nand2_1 U18768 ( .ip1(n19170), .ip2(n17082), .op(n20866) );
  inv_1 U18769 ( .ip(n20866), .op(n17086) );
  inv_1 U18770 ( .ip(n20871), .op(n17084) );
  nor2_1 U18771 ( .ip1(n17083), .ip2(n19172), .op(n20869) );
  nand2_1 U18772 ( .ip1(n17084), .ip2(n20869), .op(n17085) );
  nor2_1 U18773 ( .ip1(n20865), .ip2(n17087), .op(n17088) );
  nor2_1 U18774 ( .ip1(n20861), .ip2(n17088), .op(n17093) );
  inv_1 U18775 ( .ip(n20869), .op(n17089) );
  nor2_1 U18776 ( .ip1(n20876), .ip2(n17089), .op(n19042) );
  inv_1 U18777 ( .ip(n20865), .op(n17090) );
  nand2_1 U18778 ( .ip1(n19042), .ip2(n17090), .op(n17091) );
  or2_1 U18779 ( .ip1(n17091), .ip2(n19177), .op(n17092) );
  nand2_1 U18780 ( .ip1(n17093), .ip2(n17092), .op(n17094) );
  xnor2_1 U18781 ( .ip1(n17095), .ip2(n17094), .op(n17096) );
  nand2_1 U18782 ( .ip1(n17096), .ip2(n21577), .op(n17127) );
  and2_1 U18783 ( .ip1(n19427), .ip2(n17097), .op(n17098) );
  and2_1 U18784 ( .ip1(n17121), .ip2(n17098), .op(n17140) );
  nand2_1 U18785 ( .ip1(n17099), .ip2(n20911), .op(n17105) );
  nand2_1 U18786 ( .ip1(n10181), .ip2(n17100), .op(n17101) );
  nand2_1 U18787 ( .ip1(n17101), .ip2(n21557), .op(n17104) );
  nand3_1 U18788 ( .ip1(n17073), .ip2(n20904), .ip3(n17102), .op(n17103) );
  nand4_1 U18789 ( .ip1(n17105), .ip2(n20735), .ip3(n17104), .ip4(n17103), 
        .op(n17117) );
  nor2_1 U18790 ( .ip1(n18936), .ip2(n17167), .op(n17114) );
  nand2_1 U18791 ( .ip1(n17106), .ip2(n21540), .op(n17112) );
  nor2_1 U18792 ( .ip1(n10191), .ip2(n17269), .op(n17107) );
  not_ab_or_c_or_d U18793 ( .ip1(n21536), .ip2(n19068), .ip3(n18918), .ip4(
        n17107), .op(n17110) );
  nand2_1 U18794 ( .ip1(n18927), .ip2(n17073), .op(n17109) );
  nand2_1 U18795 ( .ip1(n19056), .ip2(n19199), .op(n17108) );
  nand3_1 U18796 ( .ip1(n17110), .ip2(n17109), .ip3(n17108), .op(n17111) );
  nand3_1 U18797 ( .ip1(n17112), .ip2(n20900), .ip3(n17111), .op(n17113) );
  not_ab_or_c_or_d U18798 ( .ip1(n17115), .ip2(n19193), .ip3(n17114), .ip4(
        n17113), .op(n17116) );
  not_ab_or_c_or_d U18799 ( .ip1(n17523), .ip2(n17140), .ip3(n17117), .ip4(
        n17116), .op(n17126) );
  nor2_1 U18800 ( .ip1(n20887), .ip2(n17178), .op(n17119) );
  nor2_1 U18801 ( .ip1(n13881), .ip2(n17184), .op(n17118) );
  not_ab_or_c_or_d U18802 ( .ip1(n17120), .ip2(n19427), .ip3(n17119), .ip4(
        n17118), .op(n17153) );
  nand2_1 U18803 ( .ip1(n17153), .ip2(n19213), .op(n17125) );
  nand2_1 U18804 ( .ip1(n17121), .ip2(n18913), .op(n17122) );
  mux2_1 U18805 ( .ip1(n20905), .ip2(n17122), .s(n19427), .op(n17123) );
  nand2_1 U18806 ( .ip1(n17123), .ip2(n18916), .op(n17154) );
  nand2_1 U18807 ( .ip1(n17154), .ip2(n19205), .op(n17124) );
  nand2_1 U18808 ( .ip1(n17129), .ip2(n17128), .op(n17138) );
  inv_1 U18809 ( .ip(n17130), .op(n20212) );
  nor2_1 U18810 ( .ip1(n17133), .ip2(n20212), .op(n17131) );
  nor2_1 U18811 ( .ip1(n17132), .ip2(n17131), .op(n17136) );
  inv_1 U18812 ( .ip(n17133), .op(n20208) );
  nand2_1 U18813 ( .ip1(n20209), .ip2(n20208), .op(n17134) );
  or2_1 U18814 ( .ip1(n17134), .ip2(n20717), .op(n17135) );
  nand2_1 U18815 ( .ip1(n17136), .ip2(n17135), .op(n17137) );
  xnor2_1 U18816 ( .ip1(n17138), .ip2(n17137), .op(n17139) );
  nand2_1 U18817 ( .ip1(n17139), .ip2(n21577), .op(n17158) );
  nand2_1 U18818 ( .ip1(n17140), .ip2(n19429), .op(n17148) );
  nand2_1 U18819 ( .ip1(n17141), .ip2(n20911), .op(n17147) );
  nand3_1 U18820 ( .ip1(n17142), .ip2(n20904), .ip3(n12138), .op(n17146) );
  nand2_1 U18821 ( .ip1(n16506), .ip2(n17143), .op(n17144) );
  nand2_1 U18822 ( .ip1(n17144), .ip2(n21557), .op(n17145) );
  nor2_1 U18823 ( .ip1(n20726), .ip2(n17149), .op(n17150) );
  not_ab_or_c_or_d U18824 ( .ip1(n20736), .ip2(n17152), .ip3(n17151), .ip4(
        n17150), .op(n17157) );
  nand2_1 U18825 ( .ip1(n17153), .ip2(n20900), .op(n17156) );
  nand2_1 U18826 ( .ip1(n17154), .ip2(n20239), .op(n17155) );
  nand2_1 U18827 ( .ip1(n17160), .ip2(n17159), .op(n17164) );
  or2_1 U18828 ( .ip1(n17161), .ip2(n19177), .op(n17162) );
  nand2_1 U18829 ( .ip1(n17515), .ip2(n17162), .op(n17163) );
  xnor2_1 U18830 ( .ip1(n17164), .ip2(n17163), .op(n17165) );
  nand2_1 U18831 ( .ip1(n17165), .ip2(n21577), .op(n17190) );
  nand2_1 U18832 ( .ip1(n17166), .ip2(n17529), .op(n17169) );
  nand2_1 U18833 ( .ip1(n17167), .ip2(n17541), .op(n17168) );
  nand2_1 U18834 ( .ip1(n17169), .ip2(n17168), .op(n17183) );
  nand2_1 U18835 ( .ip1(n17170), .ip2(n18367), .op(n17181) );
  nand2_1 U18836 ( .ip1(n10849), .ip2(n17171), .op(n17172) );
  nand2_1 U18837 ( .ip1(n17172), .ip2(n21557), .op(n17175) );
  nand3_1 U18838 ( .ip1(n18737), .ip2(n20904), .ip3(n17173), .op(n17174) );
  nand2_1 U18839 ( .ip1(n17175), .ip2(n17174), .op(n17176) );
  not_ab_or_c_or_d U18840 ( .ip1(n20911), .ip2(n17177), .ip3(n19066), .ip4(
        n17176), .op(n17180) );
  nand2_1 U18841 ( .ip1(n17178), .ip2(n18374), .op(n17179) );
  nand3_1 U18842 ( .ip1(n17181), .ip2(n17180), .ip3(n17179), .op(n17182) );
  not_ab_or_c_or_d U18843 ( .ip1(n17547), .ip2(n17184), .ip3(n17183), .ip4(
        n17182), .op(n17189) );
  nand2_1 U18844 ( .ip1(n17185), .ip2(n19205), .op(n17188) );
  nand2_1 U18845 ( .ip1(n17186), .ip2(n17523), .op(n17187) );
  nand2_1 U18846 ( .ip1(n17192), .ip2(n17191), .op(n17197) );
  nor2_1 U18847 ( .ip1(n17193), .ip2(n17565), .op(n17195) );
  nor2_1 U18848 ( .ip1(n17195), .ip2(n17194), .op(n17196) );
  nand2_1 U18849 ( .ip1(n17198), .ip2(n21577), .op(n17242) );
  inv_1 U18850 ( .ip(n20911), .op(n21555) );
  nor2_1 U18851 ( .ip1(n21555), .ip2(n10177), .op(n17221) );
  nor2_1 U18852 ( .ip1(n17199), .ip2(n10185), .op(n17200) );
  nor2_1 U18853 ( .ip1(n20907), .ip2(n17200), .op(n17220) );
  and3_1 U18854 ( .ip1(n10185), .ip2(n20904), .ip3(n17199), .op(n17219) );
  inv_1 U18855 ( .ip(n17201), .op(n17202) );
  nor2_1 U18856 ( .ip1(n20887), .ip2(n17202), .op(n17217) );
  nand2_1 U18857 ( .ip1(n21536), .ip2(n12932), .op(n17206) );
  nand2_1 U18858 ( .ip1(n18927), .ip2(n10185), .op(n17205) );
  nand2_1 U18859 ( .ip1(n20892), .ip2(n10187), .op(n17204) );
  nand2_1 U18860 ( .ip1(n19056), .ip2(n13022), .op(n17203) );
  nor2_1 U18861 ( .ip1(n18918), .ip2(n21541), .op(n17216) );
  nor2_1 U18862 ( .ip1(n17227), .ip2(n17207), .op(n17214) );
  nor2_1 U18863 ( .ip1(n17237), .ip2(n17208), .op(n17213) );
  nor2_1 U18864 ( .ip1(n17223), .ip2(n17209), .op(n17212) );
  nor2_1 U18865 ( .ip1(n17443), .ip2(n17210), .op(n17211) );
  nor2_1 U18866 ( .ip1(n20736), .ip2(n20737), .op(n17215) );
  nor2_1 U18867 ( .ip1(n17223), .ip2(n17222), .op(n17231) );
  nor2_1 U18868 ( .ip1(n17237), .ip2(n17224), .op(n17230) );
  nor2_1 U18869 ( .ip1(n17443), .ip2(n17225), .op(n17229) );
  nor2_1 U18870 ( .ip1(n17227), .ip2(n17226), .op(n17228) );
  or4_1 U18871 ( .ip1(n17231), .ip2(n17230), .ip3(n17229), .ip4(n17228), .op(
        n20725) );
  inv_1 U18872 ( .ip(n20725), .op(n17232) );
  mux2_1 U18873 ( .ip1(n20733), .ip2(n17232), .s(n13881), .op(n17233) );
  nand2_1 U18874 ( .ip1(n17233), .ip2(n21544), .op(n17234) );
  mux2_1 U18875 ( .ip1(n20735), .ip2(n17234), .s(n20885), .op(n17240) );
  mux2_1 U18876 ( .ip1(n17236), .ip2(n17235), .s(n17575), .op(n17238) );
  and2_1 U18877 ( .ip1(n17238), .ip2(n17237), .op(n19047) );
  nand2_1 U18878 ( .ip1(n19047), .ip2(n21562), .op(n17239) );
  nand2_1 U18879 ( .ip1(n17244), .ip2(n17243), .op(n17265) );
  inv_1 U18880 ( .ip(n17245), .op(n17249) );
  nor2_1 U18881 ( .ip1(n17247), .ip2(n17246), .op(n17248) );
  nor2_1 U18882 ( .ip1(n17249), .ip2(n17248), .op(n17254) );
  nand2_1 U18883 ( .ip1(n17251), .ip2(n17250), .op(n17256) );
  or2_1 U18884 ( .ip1(n17256), .ip2(n17252), .op(n17253) );
  nand2_1 U18885 ( .ip1(n17254), .ip2(n17253), .op(n17259) );
  nor2_1 U18886 ( .ip1(n17256), .ip2(n17255), .op(n17260) );
  and2_1 U18887 ( .ip1(n17260), .ip2(n17257), .op(n17258) );
  nor2_1 U18888 ( .ip1(n17259), .ip2(n17258), .op(n17263) );
  nand2_1 U18889 ( .ip1(n17260), .ip2(n19417), .op(n17261) );
  or2_1 U18890 ( .ip1(n17261), .ip2(n20717), .op(n17262) );
  nand2_1 U18891 ( .ip1(n17263), .ip2(n17262), .op(n17264) );
  xnor2_1 U18892 ( .ip1(n17265), .ip2(n17264), .op(n17266) );
  nand2_1 U18893 ( .ip1(n17266), .ip2(n21577), .op(n17295) );
  inv_1 U18894 ( .ip(n19050), .op(n17287) );
  nor2_1 U18895 ( .ip1(n17267), .ip2(n16526), .op(n17274) );
  nor2_1 U18896 ( .ip1(n10190), .ip2(n17268), .op(n17273) );
  nor2_1 U18897 ( .ip1(n10517), .ip2(n17269), .op(n17272) );
  nor2_1 U18898 ( .ip1(n11180), .ip2(n21532), .op(n17271) );
  nor2_1 U18899 ( .ip1(n17275), .ip2(n19059), .op(n17286) );
  inv_1 U18900 ( .ip(n19060), .op(n17276) );
  nand2_1 U18901 ( .ip1(n17276), .ip2(n17529), .op(n17284) );
  nand2_1 U18902 ( .ip1(n11180), .ip2(n17277), .op(n17279) );
  nor3_1 U18903 ( .ip1(n17277), .ip2(n21551), .ip3(n11180), .op(n17278) );
  not_ab_or_c_or_d U18904 ( .ip1(n21557), .ip2(n17279), .ip3(n17278), .ip4(
        n19066), .op(n17283) );
  nand2_1 U18905 ( .ip1(n19046), .ip2(n18367), .op(n17282) );
  or2_1 U18906 ( .ip1(n21555), .ip2(n17280), .op(n17281) );
  not_ab_or_c_or_d U18907 ( .ip1(n18374), .ip2(n17287), .ip3(n17286), .ip4(
        n17285), .op(n17294) );
  inv_1 U18908 ( .ip(n20733), .op(n17288) );
  nor2_1 U18909 ( .ip1(n20726), .ip2(n17288), .op(n17290) );
  nor2_1 U18910 ( .ip1(n17498), .ip2(n20725), .op(n17289) );
  nor2_1 U18911 ( .ip1(n17290), .ip2(n17289), .op(n17291) );
  mux2_1 U18912 ( .ip1(n19064), .ip2(n17291), .s(n20885), .op(n17293) );
  nand2_1 U18913 ( .ip1(n19047), .ip2(n17547), .op(n17292) );
  nand2_1 U18914 ( .ip1(n17299), .ip2(n17298), .op(n21426) );
  nor2_1 U18915 ( .ip1(n22059), .ip2(n21426), .op(n17374) );
  nor2_1 U18916 ( .ip1(n21414), .ip2(n17374), .op(n17300) );
  xor2_1 U18917 ( .ip1(n22061), .ip2(n17300), .op(n17304) );
  nor2_1 U18918 ( .ip1(n17301), .ip2(n22665), .op(n17303) );
  nor2_1 U18919 ( .ip1(n21425), .ip2(n21680), .op(n17302) );
  ab_or_c_or_d U18920 ( .ip1(n22042), .ip2(n17304), .ip3(n17303), .ip4(n17302), 
        .op(n22850) );
  nand2_1 U18921 ( .ip1(n20965), .ip2(n17305), .op(n21168) );
  inv_1 U18922 ( .ip(n21168), .op(n21043) );
  nor2_1 U18923 ( .ip1(n21043), .ip2(n10364), .op(n21174) );
  inv_1 U18924 ( .ip(\pipeline/PC_WB [8]), .op(n17308) );
  nand2_1 U18925 ( .ip1(\pipeline/PC_WB [6]), .ip2(\pipeline/PC_WB [7]), .op(
        n17307) );
  nand2_1 U18926 ( .ip1(\pipeline/PC_WB [3]), .ip2(\pipeline/PC_WB [4]), .op(
        n17306) );
  nand2_1 U18927 ( .ip1(n20972), .ip2(\pipeline/PC_WB [2]), .op(n21169) );
  nor2_1 U18928 ( .ip1(n17306), .ip2(n21169), .op(n21044) );
  nand2_1 U18929 ( .ip1(n21044), .ip2(\pipeline/PC_WB [5]), .op(n17998) );
  nor2_1 U18930 ( .ip1(n17307), .ip2(n17998), .op(n19682) );
  xor2_1 U18931 ( .ip1(n17308), .ip2(n19682), .op(n17309) );
  nand2_1 U18932 ( .ip1(n10364), .ip2(n21168), .op(n21171) );
  nor2_1 U18933 ( .ip1(n17309), .ip2(n21171), .op(n17311) );
  nor2_1 U18934 ( .ip1(n21168), .ip2(n19700), .op(n17310) );
  ab_or_c_or_d U18935 ( .ip1(n21174), .ip2(\pipeline/epc [8]), .ip3(n17311), 
        .ip4(n17310), .op(n22851) );
  inv_1 U18936 ( .ip(\pipeline/PC_WB [11]), .op(n17313) );
  nand2_1 U18937 ( .ip1(\pipeline/PC_WB [9]), .ip2(\pipeline/PC_WB [10]), .op(
        n17312) );
  nand2_1 U18938 ( .ip1(n19682), .ip2(\pipeline/PC_WB [8]), .op(n19771) );
  nor2_1 U18939 ( .ip1(n17312), .ip2(n19771), .op(n19773) );
  xor2_1 U18940 ( .ip1(n17313), .ip2(n19773), .op(n17314) );
  nor2_1 U18941 ( .ip1(n21171), .ip2(n17314), .op(n17316) );
  nor2_1 U18942 ( .ip1(n21168), .ip2(n20196), .op(n17315) );
  ab_or_c_or_d U18943 ( .ip1(n21174), .ip2(\pipeline/epc [11]), .ip3(n17316), 
        .ip4(n17315), .op(n22852) );
  nor2_1 U18944 ( .ip1(n17317), .ip2(n17628), .op(n18691) );
  inv_1 U18945 ( .ip(n18691), .op(n17318) );
  nand2_1 U18946 ( .ip1(n20965), .ip2(n22112), .op(n21210) );
  nor2_1 U18947 ( .ip1(n17318), .ip2(n21210), .op(n17323) );
  inv_1 U18948 ( .ip(\pipeline/ctrl/prev_killed_WB ), .op(n17319) );
  nand2_1 U18949 ( .ip1(n20972), .ip2(n17319), .op(n17321) );
  nor2_1 U18950 ( .ip1(n17321), .ip2(n17320), .op(n17358) );
  inv_1 U18951 ( .ip(n17358), .op(n17322) );
  nand2_1 U18952 ( .ip1(n17322), .ip2(n20966), .op(n17352) );
  nor2_1 U18953 ( .ip1(n17323), .ip2(n17352), .op(n21117) );
  inv_1 U18954 ( .ip(\pipeline/csr/instret_full [43]), .op(n17328) );
  inv_1 U18955 ( .ip(\pipeline/csr/instret_full [42]), .op(n18478) );
  inv_1 U18956 ( .ip(\pipeline/csr/instret_full [40]), .op(n18401) );
  inv_1 U18957 ( .ip(\pipeline/csr/instret_full [38]), .op(n20339) );
  inv_1 U18958 ( .ip(\pipeline/csr/instret_full [36]), .op(n20810) );
  inv_1 U18959 ( .ip(\pipeline/csr/instret_full [34]), .op(n21114) );
  inv_1 U18960 ( .ip(\pipeline/csr/instret_full [32]), .op(n20840) );
  inv_1 U18961 ( .ip(\pipeline/csr/instret_full [24]), .op(n18786) );
  inv_1 U18962 ( .ip(\pipeline/csr/instret_full [22]), .op(n20093) );
  inv_1 U18963 ( .ip(\pipeline/csr/instret_full [18]), .op(n18558) );
  inv_1 U18964 ( .ip(\pipeline/csr/instret_full [16]), .op(n19944) );
  inv_1 U18965 ( .ip(\pipeline/csr/instret_full [14]), .op(n19881) );
  inv_1 U18966 ( .ip(\pipeline/csr/instret_full [10]), .op(n19821) );
  inv_1 U18967 ( .ip(\pipeline/csr/instret_full [6]), .op(n20370) );
  nand2_1 U18968 ( .ip1(\pipeline/csr/instret_full [0]), .ip2(
        \pipeline/csr/instret_full [1]), .op(n20997) );
  nor2_1 U18969 ( .ip1(n20998), .ip2(n20997), .op(n21002) );
  nand2_1 U18970 ( .ip1(\pipeline/csr/instret_full [3]), .ip2(n21002), .op(
        n21008) );
  nor2_1 U18971 ( .ip1(n21009), .ip2(n21008), .op(n17823) );
  nand2_1 U18972 ( .ip1(\pipeline/csr/instret_full [5]), .ip2(n17823), .op(
        n20371) );
  nor2_1 U18973 ( .ip1(n20370), .ip2(n20371), .op(n20369) );
  nand2_1 U18974 ( .ip1(\pipeline/csr/instret_full [7]), .ip2(n20369), .op(
        n17367) );
  inv_1 U18975 ( .ip(\pipeline/csr/instret_full [8]), .op(n17366) );
  nor2_1 U18976 ( .ip1(n17367), .ip2(n17366), .op(n18410) );
  nand2_1 U18977 ( .ip1(\pipeline/csr/instret_full [9]), .ip2(n18410), .op(
        n19818) );
  nor2_1 U18978 ( .ip1(n19821), .ip2(n19818), .op(n17354) );
  nand2_1 U18979 ( .ip1(\pipeline/csr/instret_full [11]), .ip2(n17354), .op(
        n20780) );
  nor2_1 U18980 ( .ip1(n20781), .ip2(n20780), .op(n18051) );
  nand2_1 U18981 ( .ip1(\pipeline/csr/instret_full [13]), .ip2(n18051), .op(
        n19878) );
  nor2_1 U18982 ( .ip1(n19881), .ip2(n19878), .op(n19476) );
  nand2_1 U18983 ( .ip1(\pipeline/csr/instret_full [15]), .ip2(n19476), .op(
        n19941) );
  nor2_1 U18984 ( .ip1(n19944), .ip2(n19941), .op(n19993) );
  nand2_1 U18985 ( .ip1(\pipeline/csr/instret_full [17]), .ip2(n19993), .op(
        n18554) );
  nor2_1 U18986 ( .ip1(n18558), .ip2(n18554), .op(n18615) );
  nand2_1 U18987 ( .ip1(\pipeline/csr/instret_full [19]), .ip2(n18615), .op(
        n19540) );
  nor2_1 U18988 ( .ip1(n19541), .ip2(n19540), .op(n18679) );
  nand2_1 U18989 ( .ip1(\pipeline/csr/instret_full [21]), .ip2(n18679), .op(
        n20090) );
  nor2_1 U18990 ( .ip1(n20093), .ip2(n20090), .op(n18780) );
  nand2_1 U18991 ( .ip1(\pipeline/csr/instret_full [23]), .ip2(n18780), .op(
        n18785) );
  nor2_1 U18992 ( .ip1(n18786), .ip2(n18785), .op(n18818) );
  nand2_1 U18993 ( .ip1(\pipeline/csr/instret_full [25]), .ip2(n18818), .op(
        n19122) );
  nor2_1 U18994 ( .ip1(n19125), .ip2(n19122), .op(n19145) );
  nand2_1 U18995 ( .ip1(\pipeline/csr/instret_full [27]), .ip2(n19145), .op(
        n19284) );
  nor2_1 U18996 ( .ip1(n19287), .ip2(n19284), .op(n18892) );
  and2_1 U18997 ( .ip1(\pipeline/csr/instret_full [29]), .ip2(n18892), .op(
        n18894) );
  inv_1 U18998 ( .ip(n18894), .op(n19005) );
  nor2_1 U18999 ( .ip1(n19006), .ip2(n19005), .op(n20954) );
  nand2_1 U19000 ( .ip1(\pipeline/csr/instret_full [31]), .ip2(n20954), .op(
        n20841) );
  nor2_1 U19001 ( .ip1(n20840), .ip2(n20841), .op(n21105) );
  nand2_1 U19002 ( .ip1(\pipeline/csr/instret_full [33]), .ip2(n21105), .op(
        n21113) );
  nor2_1 U19003 ( .ip1(n21114), .ip2(n21113), .op(n21112) );
  nand2_1 U19004 ( .ip1(\pipeline/csr/instret_full [35]), .ip2(n21112), .op(
        n20811) );
  nor2_1 U19005 ( .ip1(n20810), .ip2(n20811), .op(n20809) );
  nand2_1 U19006 ( .ip1(\pipeline/csr/instret_full [37]), .ip2(n20809), .op(
        n20340) );
  nor2_1 U19007 ( .ip1(n20339), .ip2(n20340), .op(n20338) );
  nand2_1 U19008 ( .ip1(\pipeline/csr/instret_full [39]), .ip2(n20338), .op(
        n18400) );
  nor2_1 U19009 ( .ip1(n18401), .ip2(n18400), .op(n18471) );
  nand2_1 U19010 ( .ip1(\pipeline/csr/instret_full [41]), .ip2(n18471), .op(
        n18477) );
  nor2_1 U19011 ( .ip1(n18478), .ip2(n18477), .op(n18476) );
  inv_1 U19012 ( .ip(n18476), .op(n17327) );
  nand2_1 U19013 ( .ip1(\pipeline/csr/instret_full [43]), .ip2(n18476), .op(
        n18481) );
  inv_1 U19014 ( .ip(n18481), .op(n17326) );
  nor2_1 U19015 ( .ip1(htif_reset), .ip2(n21210), .op(n17361) );
  inv_1 U19016 ( .ip(n17361), .op(n17356) );
  nor2_1 U19017 ( .ip1(n18691), .ip2(n17358), .op(n17324) );
  nor2_1 U19018 ( .ip1(n17356), .ip2(n17324), .op(n18695) );
  nand2_1 U19019 ( .ip1(n17778), .ip2(n22092), .op(n17632) );
  nor2_1 U19020 ( .ip1(\pipeline/inst_DX [27]), .ip2(n17632), .op(n17360) );
  or2_1 U19021 ( .ip1(n17360), .ip2(n17632), .op(n18690) );
  nand2_1 U19022 ( .ip1(n18695), .ip2(n18690), .op(n17325) );
  inv_1 U19023 ( .ip(htif_reset), .op(n20966) );
  nand2_1 U19024 ( .ip1(n21210), .ip2(n20966), .op(n22257) );
  inv_1 U19025 ( .ip(n22257), .op(n21120) );
  buf_1 U19026 ( .ip(n21120), .op(n21217) );
  nand2_1 U19027 ( .ip1(n17358), .ip2(n21217), .op(n21010) );
  and2_1 U19028 ( .ip1(n17325), .ip2(n21010), .op(n21111) );
  not_ab_or_c_or_d U19029 ( .ip1(n17328), .ip2(n17327), .ip3(n17326), .ip4(
        n21111), .op(n17330) );
  nand2_1 U19030 ( .ip1(n17361), .ip2(n18691), .op(n21110) );
  nor2_1 U19031 ( .ip1(n21110), .ip2(n20196), .op(n17329) );
  ab_or_c_or_d U19032 ( .ip1(n21117), .ip2(\pipeline/csr/instret_full [43]), 
        .ip3(n17330), .ip4(n17329), .op(n22853) );
  fulladder U19033 ( .a(\pipeline/md/a [1]), .b(n17331), .ci(n21501), .co(
        n17340), .s(n17339) );
  inv_1 U19034 ( .ip(\pipeline/md/a [1]), .op(n17332) );
  nor2_1 U19035 ( .ip1(n17332), .ip2(n14770), .op(n17338) );
  nand2_1 U19036 ( .ip1(n21649), .ip2(n21500), .op(n17333) );
  nand2_1 U19037 ( .ip1(n20649), .ip2(n17333), .op(n17336) );
  nand2_1 U19038 ( .ip1(n21649), .ip2(n21624), .op(n20647) );
  nor2_1 U19039 ( .ip1(n21500), .ip2(n20647), .op(n17335) );
  mux2_1 U19040 ( .ip1(n17336), .ip2(n17335), .s(n17334), .op(n17337) );
  ab_or_c_or_d U19041 ( .ip1(n21944), .ip2(n17339), .ip3(n17338), .ip4(n17337), 
        .op(n22854) );
  fulladder U19042 ( .a(n17341), .b(\pipeline/md/a [2]), .ci(n17340), .co(
        n17850), .s(n17350) );
  nor2_1 U19043 ( .ip1(n17342), .ip2(n14770), .op(n17349) );
  nand2_1 U19044 ( .ip1(n21649), .ip2(n17344), .op(n17343) );
  nand2_1 U19045 ( .ip1(n20649), .ip2(n17343), .op(n17347) );
  nor2_1 U19046 ( .ip1(n17344), .ip2(n20647), .op(n17346) );
  mux2_1 U19047 ( .ip1(n17347), .ip2(n17346), .s(n17345), .op(n17348) );
  ab_or_c_or_d U19048 ( .ip1(n21944), .ip2(n17350), .ip3(n17349), .ip4(n17348), 
        .op(n22855) );
  inv_1 U19049 ( .ip(n17360), .op(n17351) );
  nor2_1 U19050 ( .ip1(n17351), .ip2(n21210), .op(n17353) );
  nor2_1 U19051 ( .ip1(n17353), .ip2(n17352), .op(n21016) );
  inv_1 U19052 ( .ip(\pipeline/csr/instret_full [11]), .op(n17355) );
  mux2_1 U19053 ( .ip1(n17355), .ip2(\pipeline/csr/instret_full [11]), .s(
        n17354), .op(n17359) );
  nor2_1 U19054 ( .ip1(n17360), .ip2(n17356), .op(n17357) );
  nand2_1 U19055 ( .ip1(n17358), .ip2(n17357), .op(n18555) );
  and2_1 U19056 ( .ip1(n21010), .ip2(n18555), .op(n21005) );
  nor2_1 U19057 ( .ip1(n17359), .ip2(n21005), .op(n17363) );
  nand2_1 U19058 ( .ip1(n17361), .ip2(n17360), .op(n21001) );
  nor2_1 U19059 ( .ip1(n21001), .ip2(n20196), .op(n17362) );
  ab_or_c_or_d U19060 ( .ip1(n21016), .ip2(\pipeline/csr/instret_full [11]), 
        .ip3(n17363), .ip4(n17362), .op(n22856) );
  nand2_1 U19061 ( .ip1(n20965), .ip2(n17364), .op(n21029) );
  nor2_1 U19062 ( .ip1(n21029), .ip2(n19700), .op(n17365) );
  ab_or_c_or_d U19063 ( .ip1(\pipeline/csr/mtvec [8]), .ip2(n21029), .ip3(
        htif_reset), .ip4(n17365), .op(n22857) );
  not_ab_or_c_or_d U19064 ( .ip1(n17367), .ip2(n17366), .ip3(n18410), .ip4(
        n21005), .op(n17369) );
  nor2_1 U19065 ( .ip1(n21001), .ip2(n19700), .op(n17368) );
  ab_or_c_or_d U19066 ( .ip1(n21016), .ip2(\pipeline/csr/instret_full [8]), 
        .ip3(n17369), .ip4(n17368), .op(n22858) );
  nor2_1 U19067 ( .ip1(n22619), .ip2(n22665), .op(n17384) );
  inv_1 U19068 ( .ip(n21360), .op(n21406) );
  or2_1 U19069 ( .ip1(n22062), .ip2(n22064), .op(n17379) );
  inv_1 U19070 ( .ip(n22065), .op(n17372) );
  inv_1 U19071 ( .ip(n17370), .op(n17371) );
  nand2_1 U19072 ( .ip1(n17372), .ip2(n17371), .op(n17375) );
  inv_1 U19073 ( .ip(n22061), .op(n17373) );
  nand2_1 U19074 ( .ip1(n17374), .ip2(n17373), .op(n21420) );
  nor2_1 U19075 ( .ip1(n17375), .ip2(n21420), .op(n21407) );
  nor2_1 U19076 ( .ip1(n17376), .ip2(n22052), .op(n17377) );
  nand2_1 U19077 ( .ip1(n21407), .ip2(n17377), .op(n21393) );
  nor2_1 U19078 ( .ip1(n22054), .ip2(n21393), .op(n17410) );
  inv_1 U19079 ( .ip(n22056), .op(n17378) );
  nand2_1 U19080 ( .ip1(n17410), .ip2(n17378), .op(n21387) );
  nor2_1 U19081 ( .ip1(n22058), .ip2(n21387), .op(n21381) );
  inv_1 U19082 ( .ip(n22060), .op(n21383) );
  nand2_1 U19083 ( .ip1(n21381), .ip2(n21383), .op(n21374) );
  nor2_1 U19084 ( .ip1(n17379), .ip2(n21374), .op(n17386) );
  nor2_1 U19085 ( .ip1(n21406), .ip2(n17386), .op(n17382) );
  nand2_1 U19086 ( .ip1(n17386), .ip2(n22042), .op(n17380) );
  nand2_1 U19087 ( .ip1(n17380), .ip2(n21409), .op(n17381) );
  mux2_1 U19088 ( .ip1(n17382), .ip2(n17381), .s(n22068), .op(n17383) );
  ab_or_c_or_d U19089 ( .ip1(n21493), .ip2(\pipeline/md/b [46]), .ip3(n17384), 
        .ip4(n17383), .op(n22859) );
  nor2_1 U19090 ( .ip1(n22680), .ip2(n22665), .op(n17396) );
  inv_1 U19091 ( .ip(n22068), .op(n17385) );
  nand2_1 U19092 ( .ip1(n17386), .ip2(n17385), .op(n21361) );
  nor2_1 U19093 ( .ip1(n22082), .ip2(n21361), .op(n21354) );
  inv_1 U19094 ( .ip(n17387), .op(n17388) );
  nand2_1 U19095 ( .ip1(n21354), .ip2(n17388), .op(n21349) );
  nor2_1 U19096 ( .ip1(n22083), .ip2(n21349), .op(n21343) );
  inv_1 U19097 ( .ip(n22084), .op(n17389) );
  nand2_1 U19098 ( .ip1(n21343), .ip2(n17389), .op(n21336) );
  nor2_1 U19099 ( .ip1(n22085), .ip2(n21336), .op(n17402) );
  nand2_1 U19100 ( .ip1(n17402), .ip2(n22042), .op(n17390) );
  nand2_1 U19101 ( .ip1(n17390), .ip2(n21409), .op(n17394) );
  nor2_1 U19102 ( .ip1(n21406), .ip2(n17402), .op(n17393) );
  nand2_1 U19103 ( .ip1(n17392), .ip2(n17391), .op(n17427) );
  mux2_1 U19104 ( .ip1(n17394), .ip2(n17393), .s(n17427), .op(n17395) );
  ab_or_c_or_d U19105 ( .ip1(n21493), .ip2(\pipeline/md/b [52]), .ip3(n17396), 
        .ip4(n17395), .op(n22860) );
  nor2_1 U19106 ( .ip1(n22699), .ip2(n22665), .op(n17409) );
  inv_1 U19107 ( .ip(n19308), .op(n17397) );
  or2_1 U19108 ( .ip1(n17397), .ip2(n17399), .op(n17401) );
  nand2_1 U19109 ( .ip1(n17399), .ip2(n17398), .op(n17400) );
  nand2_1 U19110 ( .ip1(n17401), .ip2(n17400), .op(n22086) );
  nand2_1 U19111 ( .ip1(n17402), .ip2(n17427), .op(n21331) );
  nor2_1 U19112 ( .ip1(n22086), .ip2(n21331), .op(n21280) );
  nand2_1 U19113 ( .ip1(n21280), .ip2(n22042), .op(n17403) );
  nand2_1 U19114 ( .ip1(n17403), .ip2(n21409), .op(n17407) );
  nor2_1 U19115 ( .ip1(n21406), .ip2(n21280), .op(n17406) );
  nand2_1 U19116 ( .ip1(n17405), .ip2(n17404), .op(n21279) );
  mux2_1 U19117 ( .ip1(n17407), .ip2(n17406), .s(n21279), .op(n17408) );
  ab_or_c_or_d U19118 ( .ip1(n21493), .ip2(\pipeline/md/b [54]), .ip3(n17409), 
        .ip4(n17408), .op(n22861) );
  nor2_1 U19119 ( .ip1(n21763), .ip2(n21680), .op(n17415) );
  nor2_1 U19120 ( .ip1(n21406), .ip2(n17410), .op(n17413) );
  nand2_1 U19121 ( .ip1(n17410), .ip2(n22042), .op(n17411) );
  nand2_1 U19122 ( .ip1(n17411), .ip2(n21409), .op(n17412) );
  mux2_1 U19123 ( .ip1(n17413), .ip2(n17412), .s(n22056), .op(n17414) );
  ab_or_c_or_d U19124 ( .ip1(n14765), .ip2(\pipeline/md/b [42]), .ip3(n17415), 
        .ip4(n17414), .op(n22862) );
  nor2_1 U19125 ( .ip1(n21168), .ip2(n22229), .op(n17426) );
  inv_1 U19126 ( .ip(\pipeline/PC_WB [28]), .op(n17424) );
  nand2_1 U19127 ( .ip1(\pipeline/PC_WB [24]), .ip2(\pipeline/PC_WB [25]), 
        .op(n17420) );
  nand2_1 U19128 ( .ip1(\pipeline/PC_WB [21]), .ip2(\pipeline/PC_WB [22]), 
        .op(n17419) );
  nand2_1 U19129 ( .ip1(\pipeline/PC_WB [18]), .ip2(\pipeline/PC_WB [19]), 
        .op(n17418) );
  nand2_1 U19130 ( .ip1(\pipeline/PC_WB [15]), .ip2(\pipeline/PC_WB [16]), 
        .op(n17417) );
  nand2_1 U19131 ( .ip1(\pipeline/PC_WB [12]), .ip2(\pipeline/PC_WB [13]), 
        .op(n17416) );
  nand2_1 U19132 ( .ip1(n19773), .ip2(\pipeline/PC_WB [11]), .op(n20699) );
  nor2_1 U19133 ( .ip1(n17416), .ip2(n20699), .op(n19839) );
  nand2_1 U19134 ( .ip1(n19839), .ip2(\pipeline/PC_WB [14]), .op(n18272) );
  nor2_1 U19135 ( .ip1(n17417), .ip2(n18272), .op(n19961) );
  nand2_1 U19136 ( .ip1(n19961), .ip2(\pipeline/PC_WB [17]), .op(n20028) );
  nor2_1 U19137 ( .ip1(n17418), .ip2(n20028), .op(n20030) );
  nand2_1 U19138 ( .ip1(n20030), .ip2(\pipeline/PC_WB [20]), .op(n20051) );
  nor2_1 U19139 ( .ip1(n17419), .ip2(n20051), .op(n20110) );
  nand2_1 U19140 ( .ip1(n20110), .ip2(\pipeline/PC_WB [23]), .op(n18827) );
  nor2_1 U19141 ( .ip1(n17420), .ip2(n18827), .op(n19080) );
  nand2_1 U19142 ( .ip1(n19080), .ip2(\pipeline/PC_WB [26]), .op(n17421) );
  inv_1 U19143 ( .ip(n17421), .op(n19150) );
  nand2_1 U19144 ( .ip1(n19150), .ip2(\pipeline/PC_WB [27]), .op(n17423) );
  nand2_1 U19145 ( .ip1(\pipeline/PC_WB [27]), .ip2(\pipeline/PC_WB [28]), 
        .op(n17422) );
  nor2_1 U19146 ( .ip1(n17422), .ip2(n17421), .op(n20320) );
  not_ab_or_c_or_d U19147 ( .ip1(n17424), .ip2(n17423), .ip3(n20320), .ip4(
        n21171), .op(n17425) );
  ab_or_c_or_d U19148 ( .ip1(n21174), .ip2(\pipeline/epc [28]), .ip3(n17426), 
        .ip4(n17425), .op(n22863) );
  inv_1 U19149 ( .ip(n17427), .op(n17428) );
  nand2_1 U19150 ( .ip1(n17741), .ip2(n20966), .op(n21582) );
  inv_1 U19151 ( .ip(n21582), .op(n22067) );
  mux2_1 U19152 ( .ip1(\pipeline/store_data_WB [21]), .ip2(n17428), .s(n17777), 
        .op(n8818) );
  inv_1 U19153 ( .ip(n21279), .op(n17430) );
  inv_1 U19154 ( .ip(n21582), .op(n17429) );
  buf_1 U19155 ( .ip(n17429), .op(n20389) );
  mux2_1 U19156 ( .ip1(\pipeline/store_data_WB [23]), .ip2(n17430), .s(n20389), 
        .op(n8816) );
  mux2_1 U19157 ( .ip1(dmem_hwdata[5]), .ip2(n17370), .s(n22067), .op(n8834)
         );
  inv_1 U19158 ( .ip(n17431), .op(n17432) );
  nor2_1 U19159 ( .ip1(n19894), .ip2(n17432), .op(n17434) );
  xor2_1 U19160 ( .ip1(n17434), .ip2(n17433), .op(imem_haddr[14]) );
  xor2_1 U19161 ( .ip1(n17436), .ip2(n17435), .op(n17438) );
  inv_1 U19162 ( .ip(n17437), .op(n21994) );
  nand2_1 U19163 ( .ip1(n17439), .ip2(n20239), .op(n17442) );
  nand2_1 U19164 ( .ip1(n17440), .ip2(n19429), .op(n17441) );
  nand2_1 U19165 ( .ip1(n17442), .ip2(n17441), .op(n17512) );
  nand2_1 U19166 ( .ip1(n17512), .ip2(n13881), .op(n17475) );
  nor2_1 U19167 ( .ip1(n17443), .ip2(n17478), .op(n17444) );
  nor2_1 U19168 ( .ip1(n13881), .ip2(n17444), .op(n17446) );
  nor2_1 U19169 ( .ip1(n20887), .ip2(n17542), .op(n17445) );
  ab_or_c_or_d U19170 ( .ip1(n19427), .ip2(n18948), .ip3(n17446), .ip4(n17445), 
        .op(n18378) );
  nor2_1 U19171 ( .ip1(n20724), .ip2(n18378), .op(n17466) );
  nand2_1 U19172 ( .ip1(n21536), .ip2(n13552), .op(n17449) );
  nand2_1 U19173 ( .ip1(n20892), .ip2(n13877), .op(n17448) );
  nand2_1 U19174 ( .ip1(n10189), .ip2(n19056), .op(n17447) );
  and4_1 U19175 ( .ip1(n17450), .ip2(n17449), .ip3(n17448), .ip4(n17447), .op(
        n17578) );
  nand2_1 U19176 ( .ip1(n21536), .ip2(n13636), .op(n17454) );
  nand2_1 U19177 ( .ip1(n13678), .ip2(n18927), .op(n17453) );
  nand2_1 U19178 ( .ip1(n20892), .ip2(n16506), .op(n17452) );
  nand2_1 U19179 ( .ip1(n13868), .ip2(n19056), .op(n17451) );
  inv_1 U19180 ( .ip(n20219), .op(n17576) );
  mux2_1 U19181 ( .ip1(n17578), .ip2(n17576), .s(n10198), .op(n17502) );
  nand2_1 U19182 ( .ip1(n17502), .ip2(n20736), .op(n17464) );
  nor3_1 U19183 ( .ip1(n17455), .ip2(n21551), .ip3(n10206), .op(n17460) );
  nor2_1 U19184 ( .ip1(n17457), .ip2(n17456), .op(n17458) );
  nor2_1 U19185 ( .ip1(n20907), .ip2(n17458), .op(n17459) );
  not_ab_or_c_or_d U19186 ( .ip1(n20911), .ip2(n17461), .ip3(n17460), .ip4(
        n17459), .op(n17463) );
  nand3_1 U19187 ( .ip1(n17464), .ip2(n17463), .ip3(n17462), .op(n17465) );
  not_ab_or_c_or_d U19188 ( .ip1(n21549), .ip2(n17467), .ip3(n17466), .ip4(
        n17465), .op(n17474) );
  xnor2_1 U19189 ( .ip1(n17470), .ip2(n20210), .op(n17471) );
  inv_1 U19190 ( .ip(n17471), .op(n17472) );
  nand2_1 U19191 ( .ip1(n21577), .ip2(n17472), .op(n17473) );
  nand3_1 U19192 ( .ip1(n17475), .ip2(n17474), .ip3(n17473), .op(dmem_haddr[9]) );
  nand2_1 U19193 ( .ip1(n17520), .ip2(n21540), .op(n17477) );
  nand2_1 U19194 ( .ip1(n20230), .ip2(n19427), .op(n17476) );
  nand2_1 U19195 ( .ip1(n17477), .ip2(n17476), .op(n17501) );
  inv_1 U19196 ( .ip(n17478), .op(n17544) );
  nand3_1 U19197 ( .ip1(n18913), .ip2(n17544), .ip3(n21562), .op(n17485) );
  and3_1 U19198 ( .ip1(n17479), .ip2(n20904), .ip3(n13525), .op(n17482) );
  or2_1 U19199 ( .ip1(n17480), .ip2(n17479), .op(n21533) );
  and2_1 U19200 ( .ip1(n21533), .ip2(n21557), .op(n17481) );
  not_ab_or_c_or_d U19201 ( .ip1(n20911), .ip2(n17483), .ip3(n17482), .ip4(
        n17481), .op(n17484) );
  nand2_1 U19202 ( .ip1(n17485), .ip2(n17484), .op(n17500) );
  inv_1 U19203 ( .ip(n17486), .op(n17490) );
  nand2_1 U19204 ( .ip1(n21536), .ip2(n13022), .op(n17487) );
  nand4_1 U19205 ( .ip1(n17490), .ip2(n17489), .ip3(n17488), .ip4(n17487), 
        .op(n17579) );
  mux2_1 U19206 ( .ip1(n17479), .ip2(n10184), .s(n21552), .op(n17491) );
  and2_1 U19207 ( .ip1(n17491), .ip2(n18913), .op(n17496) );
  mux2_1 U19208 ( .ip1(n17492), .ip2(n10185), .s(n21552), .op(n17494) );
  and2_1 U19209 ( .ip1(n17494), .ip2(n17493), .op(n17495) );
  not_ab_or_c_or_d U19210 ( .ip1(n10198), .ip2(n17579), .ip3(n17496), .ip4(
        n17495), .op(n17497) );
  nor2_1 U19211 ( .ip1(n17498), .ip2(n17497), .op(n17499) );
  not_ab_or_c_or_d U19212 ( .ip1(n21544), .ip2(n17501), .ip3(n17500), .ip4(
        n17499), .op(n17511) );
  nand2_1 U19213 ( .ip1(n17502), .ip2(n21549), .op(n17510) );
  inv_1 U19214 ( .ip(n17503), .op(n17507) );
  nand2_1 U19215 ( .ip1(n17505), .ip2(n17504), .op(n17506) );
  xor2_1 U19216 ( .ip1(n17507), .ip2(n17506), .op(n17508) );
  nand2_1 U19217 ( .ip1(n17508), .ip2(n21577), .op(n17509) );
  and3_1 U19218 ( .ip1(n17511), .ip2(n17510), .ip3(n17509), .op(n17514) );
  nand2_1 U19219 ( .ip1(n17512), .ip2(n19185), .op(n17513) );
  nand2_1 U19220 ( .ip1(n17514), .ip2(n17513), .op(dmem_haddr[1]) );
  inv_1 U19221 ( .ip(n21577), .op(n17518) );
  nand2_1 U19222 ( .ip1(n17516), .ip2(n17515), .op(n17517) );
  mux2_1 U19223 ( .ip1(n17520), .ip2(n17519), .s(n10198), .op(n20216) );
  nand2_1 U19224 ( .ip1(n20216), .ip2(n13881), .op(n17522) );
  nand2_1 U19225 ( .ip1(n20229), .ip2(n20896), .op(n17521) );
  nand2_1 U19226 ( .ip1(n17522), .ip2(n17521), .op(n17589) );
  nand2_1 U19227 ( .ip1(n17589), .ip2(n17523), .op(n17550) );
  nand4_1 U19228 ( .ip1(n17527), .ip2(n17526), .ip3(n17525), .ip4(n17524), 
        .op(n18935) );
  nor2_1 U19229 ( .ip1(n18948), .ip2(n17528), .op(n17540) );
  nand2_1 U19230 ( .ip1(n18934), .ip2(n17529), .op(n17538) );
  nand2_1 U19231 ( .ip1(n10192), .ip2(n17531), .op(n17533) );
  nor3_1 U19232 ( .ip1(n17531), .ip2(n21551), .ip3(n10192), .op(n17532) );
  not_ab_or_c_or_d U19233 ( .ip1(n21557), .ip2(n17533), .ip3(n17532), .ip4(
        n19066), .op(n17537) );
  nand2_1 U19234 ( .ip1(n18944), .ip2(n18367), .op(n17536) );
  nand2_1 U19235 ( .ip1(n17534), .ip2(n20911), .op(n17535) );
  not_ab_or_c_or_d U19236 ( .ip1(n17541), .ip2(n18935), .ip3(n17540), .ip4(
        n17539), .op(n17549) );
  nand2_1 U19237 ( .ip1(n17542), .ip2(n17575), .op(n17546) );
  nand2_1 U19238 ( .ip1(n17544), .ip2(n17543), .op(n17545) );
  nand2_1 U19239 ( .ip1(n17546), .ip2(n17545), .op(n18945) );
  nand2_1 U19240 ( .ip1(n18945), .ip2(n17547), .op(n17548) );
  nand3_1 U19241 ( .ip1(n17550), .ip2(n17549), .ip3(n17548), .op(n17551) );
  nor2_1 U19242 ( .ip1(n17552), .ip2(n17551), .op(n17560) );
  inv_1 U19243 ( .ip(n18914), .op(n17553) );
  nor2_1 U19244 ( .ip1(n17554), .ip2(n17553), .op(n17557) );
  inv_1 U19245 ( .ip(n18916), .op(n17555) );
  mux2_1 U19246 ( .ip1(n17555), .ip2(n20216), .s(n13881), .op(n17556) );
  nor2_1 U19247 ( .ip1(n17557), .ip2(n17556), .op(n17572) );
  or2_1 U19248 ( .ip1(n17558), .ip2(n17572), .op(n17559) );
  nand2_1 U19249 ( .ip1(n17560), .ip2(n17559), .op(dmem_haddr[21]) );
  inv_1 U19250 ( .ip(n17561), .op(n17563) );
  nand2_1 U19251 ( .ip1(n17563), .ip2(n17562), .op(n17569) );
  nor2_1 U19252 ( .ip1(n17565), .ip2(n17564), .op(n17566) );
  nor2_1 U19253 ( .ip1(n17567), .ip2(n17566), .op(n17568) );
  xor2_1 U19254 ( .ip1(n17569), .ip2(n17568), .op(n17570) );
  nor2_1 U19255 ( .ip1(n17573), .ip2(n17572), .op(n17574) );
  nor2_1 U19256 ( .ip1(n17571), .ip2(n17574), .op(n17595) );
  mux2_1 U19257 ( .ip1(n20230), .ip2(n17576), .s(n17575), .op(n17577) );
  nor2_1 U19258 ( .ip1(n20736), .ip2(n17577), .op(n17582) );
  nor2_1 U19259 ( .ip1(n20887), .ip2(n17578), .op(n17581) );
  nor2_1 U19260 ( .ip1(n18918), .ip2(n17579), .op(n17580) );
  or4_1 U19261 ( .ip1(n17583), .ip2(n17582), .ip3(n17581), .ip4(n17580), .op(
        n17593) );
  nor2_1 U19262 ( .ip1(n17584), .ip2(n10187), .op(n17585) );
  nor2_1 U19263 ( .ip1(n20907), .ip2(n17585), .op(n17587) );
  nor3_1 U19264 ( .ip1(n10194), .ip2(n21551), .ip3(n16446), .op(n17586) );
  not_ab_or_c_or_d U19265 ( .ip1(n20911), .ip2(n17588), .ip3(n17587), .ip4(
        n17586), .op(n17592) );
  nand2_1 U19266 ( .ip1(n17589), .ip2(n19429), .op(n17591) );
  nand2_1 U19267 ( .ip1(n18945), .ip2(n21562), .op(n17590) );
  and4_1 U19268 ( .ip1(n17593), .ip2(n17592), .ip3(n17591), .ip4(n17590), .op(
        n17594) );
  nand2_1 U19269 ( .ip1(n17595), .ip2(n17594), .op(dmem_haddr[5]) );
  nor2_1 U19270 ( .ip1(n22094), .ip2(n17628), .op(n17614) );
  inv_1 U19271 ( .ip(n17614), .op(n17596) );
  nand3_1 U19272 ( .ip1(n20966), .ip2(n17597), .ip3(n17596), .op(n18328) );
  inv_1 U19273 ( .ip(n18328), .op(n17598) );
  nor2_1 U19274 ( .ip1(htif_reset), .ip2(n17597), .op(n21179) );
  or2_1 U19275 ( .ip1(n21179), .ip2(n21120), .op(n20181) );
  nor2_1 U19276 ( .ip1(n17598), .ip2(n20181), .op(n22308) );
  inv_1 U19277 ( .ip(\pipeline/csr/cycle_full [61]), .op(n18972) );
  inv_1 U19278 ( .ip(\pipeline/csr/cycle_full [59]), .op(n19235) );
  inv_1 U19279 ( .ip(\pipeline/csr/cycle_full [57]), .op(n22310) );
  inv_1 U19280 ( .ip(\pipeline/csr/cycle_full [55]), .op(n22302) );
  inv_1 U19281 ( .ip(\pipeline/csr/cycle_full [53]), .op(n18687) );
  inv_1 U19282 ( .ip(\pipeline/csr/cycle_full [51]), .op(n18622) );
  inv_1 U19283 ( .ip(\pipeline/csr/cycle_full [49]), .op(n20000) );
  inv_1 U19284 ( .ip(\pipeline/csr/cycle_full [47]), .op(n19484) );
  inv_1 U19285 ( .ip(\pipeline/csr/cycle_full [45]), .op(n20272) );
  inv_1 U19286 ( .ip(\pipeline/csr/cycle_full [43]), .op(n20197) );
  inv_1 U19287 ( .ip(\pipeline/csr/cycle_full [41]), .op(n18467) );
  inv_1 U19288 ( .ip(\pipeline/csr/cycle_full [39]), .op(n19596) );
  inv_1 U19289 ( .ip(\pipeline/csr/cycle_full [37]), .op(n21069) );
  inv_1 U19290 ( .ip(\pipeline/csr/cycle_full [35]), .op(n21227) );
  inv_1 U19291 ( .ip(\pipeline/csr/cycle_full [33]), .op(n22030) );
  inv_1 U19292 ( .ip(\pipeline/csr/cycle_full [31]), .op(n17613) );
  inv_1 U19293 ( .ip(\pipeline/csr/cycle_full [29]), .op(n17612) );
  inv_1 U19294 ( .ip(\pipeline/csr/cycle_full [27]), .op(n17611) );
  inv_1 U19295 ( .ip(\pipeline/csr/cycle_full [25]), .op(n17610) );
  inv_1 U19296 ( .ip(\pipeline/csr/cycle_full [23]), .op(n17609) );
  inv_1 U19297 ( .ip(\pipeline/csr/cycle_full [21]), .op(n17608) );
  inv_1 U19298 ( .ip(\pipeline/csr/cycle_full [19]), .op(n17607) );
  inv_1 U19299 ( .ip(\pipeline/csr/cycle_full [17]), .op(n17606) );
  inv_1 U19300 ( .ip(\pipeline/csr/cycle_full [15]), .op(n17605) );
  inv_1 U19301 ( .ip(\pipeline/csr/cycle_full [13]), .op(n17604) );
  inv_1 U19302 ( .ip(\pipeline/csr/cycle_full [11]), .op(n17603) );
  inv_1 U19303 ( .ip(\pipeline/csr/cycle_full [9]), .op(n17602) );
  inv_1 U19304 ( .ip(\pipeline/csr/cycle_full [7]), .op(n17601) );
  inv_1 U19305 ( .ip(\pipeline/csr/cycle_full [5]), .op(n17600) );
  inv_1 U19306 ( .ip(\pipeline/csr/cycle_full [3]), .op(n17599) );
  nand3_1 U19307 ( .ip1(\pipeline/csr/cycle_full [2]), .ip2(
        \pipeline/csr/cycle_full [1]), .ip3(\pipeline/csr/cycle_full [0]), 
        .op(n21213) );
  nor2_1 U19308 ( .ip1(n17599), .ip2(n21213), .op(n21218) );
  nand2_1 U19309 ( .ip1(\pipeline/csr/cycle_full [4]), .ip2(n21218), .op(
        n21073) );
  nor2_1 U19310 ( .ip1(n17600), .ip2(n21073), .op(n21077) );
  nand2_1 U19311 ( .ip1(\pipeline/csr/cycle_full [6]), .ip2(n21077), .op(
        n20365) );
  nor2_1 U19312 ( .ip1(n17601), .ip2(n20365), .op(n19729) );
  nand2_1 U19313 ( .ip1(\pipeline/csr/cycle_full [8]), .ip2(n19729), .op(
        n19731) );
  nor2_1 U19314 ( .ip1(n17602), .ip2(n19731), .op(n19811) );
  nand2_1 U19315 ( .ip1(\pipeline/csr/cycle_full [10]), .ip2(n19811), .op(
        n20187) );
  nor2_1 U19316 ( .ip1(n17603), .ip2(n20187), .op(n20772) );
  nand2_1 U19317 ( .ip1(\pipeline/csr/cycle_full [12]), .ip2(n20772), .op(
        n20774) );
  nor2_1 U19318 ( .ip1(n17604), .ip2(n20774), .op(n20263) );
  nand2_1 U19319 ( .ip1(\pipeline/csr/cycle_full [14]), .ip2(n20263), .op(
        n19872) );
  nor2_1 U19320 ( .ip1(n17605), .ip2(n19872), .op(n19934) );
  nand2_1 U19321 ( .ip1(\pipeline/csr/cycle_full [16]), .ip2(n19934), .op(
        n19985) );
  nor2_1 U19322 ( .ip1(n17606), .ip2(n19985), .op(n19988) );
  nand2_1 U19323 ( .ip1(\pipeline/csr/cycle_full [18]), .ip2(n19988), .op(
        n18606) );
  nor2_1 U19324 ( .ip1(n17607), .ip2(n18606), .op(n19532) );
  nand2_1 U19325 ( .ip1(\pipeline/csr/cycle_full [20]), .ip2(n19532), .op(
        n19534) );
  nor2_1 U19326 ( .ip1(n17608), .ip2(n19534), .op(n20083) );
  nand2_1 U19327 ( .ip1(\pipeline/csr/cycle_full [22]), .ip2(n20083), .op(
        n20133) );
  nor2_1 U19328 ( .ip1(n17609), .ip2(n20133), .op(n20136) );
  nand2_1 U19329 ( .ip1(\pipeline/csr/cycle_full [24]), .ip2(n20136), .op(
        n18811) );
  nor2_1 U19330 ( .ip1(n17610), .ip2(n18811), .op(n19115) );
  nand2_1 U19331 ( .ip1(\pipeline/csr/cycle_full [26]), .ip2(n19115), .op(
        n19223) );
  nor2_1 U19332 ( .ip1(n17611), .ip2(n19223), .op(n19276) );
  nand2_1 U19333 ( .ip1(\pipeline/csr/cycle_full [28]), .ip2(n19276), .op(
        n19278) );
  nor2_1 U19334 ( .ip1(n17612), .ip2(n19278), .op(n18998) );
  nand2_1 U19335 ( .ip1(\pipeline/csr/cycle_full [30]), .ip2(n18998), .op(
        n20945) );
  nor2_1 U19336 ( .ip1(n17613), .ip2(n20945), .op(n22289) );
  nand2_1 U19337 ( .ip1(\pipeline/csr/cycle_full [32]), .ip2(n22289), .op(
        n22291) );
  nor2_1 U19338 ( .ip1(n22030), .ip2(n22291), .op(n22294) );
  nand2_1 U19339 ( .ip1(\pipeline/csr/cycle_full [34]), .ip2(n22294), .op(
        n22296) );
  nor2_1 U19340 ( .ip1(n21227), .ip2(n22296), .op(n21226) );
  nand2_1 U19341 ( .ip1(\pipeline/csr/cycle_full [36]), .ip2(n21226), .op(
        n21070) );
  nor2_1 U19342 ( .ip1(n21069), .ip2(n21070), .op(n21068) );
  nand2_1 U19343 ( .ip1(\pipeline/csr/cycle_full [38]), .ip2(n21068), .op(
        n20375) );
  nor2_1 U19344 ( .ip1(n19596), .ip2(n20375), .op(n19740) );
  nand2_1 U19345 ( .ip1(\pipeline/csr/cycle_full [40]), .ip2(n19740), .op(
        n19742) );
  nor2_1 U19346 ( .ip1(n18467), .ip2(n19742), .op(n19829) );
  nand2_1 U19347 ( .ip1(\pipeline/csr/cycle_full [42]), .ip2(n19829), .op(
        n20198) );
  nor2_1 U19348 ( .ip1(n20197), .ip2(n20198), .op(n20789) );
  nand2_1 U19349 ( .ip1(\pipeline/csr/cycle_full [44]), .ip2(n20789), .op(
        n20791) );
  nor2_1 U19350 ( .ip1(n20272), .ip2(n20791), .op(n20271) );
  nand2_1 U19351 ( .ip1(\pipeline/csr/cycle_full [46]), .ip2(n20271), .op(
        n19889) );
  nor2_1 U19352 ( .ip1(n19484), .ip2(n19889), .op(n19952) );
  nand2_1 U19353 ( .ip1(\pipeline/csr/cycle_full [48]), .ip2(n19952), .op(
        n20001) );
  nor2_1 U19354 ( .ip1(n20000), .ip2(n20001), .op(n19999) );
  nand2_1 U19355 ( .ip1(\pipeline/csr/cycle_full [50]), .ip2(n19999), .op(
        n18623) );
  nor2_1 U19356 ( .ip1(n18622), .ip2(n18623), .op(n19550) );
  nand2_1 U19357 ( .ip1(\pipeline/csr/cycle_full [52]), .ip2(n19550), .op(
        n19552) );
  nor2_1 U19358 ( .ip1(n18687), .ip2(n19552), .op(n20101) );
  nand2_1 U19359 ( .ip1(\pipeline/csr/cycle_full [54]), .ip2(n20101), .op(
        n22301) );
  nor2_1 U19360 ( .ip1(n22302), .ip2(n22301), .op(n22300) );
  nand2_1 U19361 ( .ip1(\pipeline/csr/cycle_full [56]), .ip2(n22300), .op(
        n22309) );
  nor2_1 U19362 ( .ip1(n22310), .ip2(n22309), .op(n22307) );
  nand2_1 U19363 ( .ip1(\pipeline/csr/cycle_full [58]), .ip2(n22307), .op(
        n19236) );
  nor2_1 U19364 ( .ip1(n19235), .ip2(n19236), .op(n19294) );
  nand2_1 U19365 ( .ip1(\pipeline/csr/cycle_full [60]), .ip2(n19294), .op(
        n19296) );
  nor2_1 U19366 ( .ip1(n18972), .ip2(n19296), .op(n22315) );
  nand2_1 U19367 ( .ip1(\pipeline/csr/cycle_full [62]), .ip2(n22315), .op(
        n22318) );
  nor2_1 U19368 ( .ip1(\pipeline/csr/cycle_full [63]), .ip2(n22318), .op(
        n17615) );
  nand2_1 U19369 ( .ip1(n17614), .ip2(n20966), .op(n18568) );
  nor2_1 U19370 ( .ip1(n18568), .ip2(n21210), .op(n22314) );
  not_ab_or_c_or_d U19371 ( .ip1(\pipeline/csr/cycle_full [63]), .ip2(n22318), 
        .ip3(n17615), .ip4(n22314), .op(n17616) );
  or2_1 U19372 ( .ip1(n22308), .ip2(n17616), .op(n17619) );
  inv_1 U19373 ( .ip(n18568), .op(n17620) );
  nand2_1 U19374 ( .ip1(n17620), .ip2(n20959), .op(n17617) );
  or2_1 U19375 ( .ip1(n17617), .ip2(n17616), .op(n17618) );
  nand2_1 U19376 ( .ip1(n17619), .ip2(n17618), .op(\pipeline/csr/N1936 ) );
  nand2_1 U19377 ( .ip1(n17620), .ip2(n22222), .op(n17625) );
  nor2_1 U19378 ( .ip1(n21210), .ip2(n17625), .op(n17623) );
  or2_1 U19379 ( .ip1(\pipeline/csr/cycle_full [58]), .ip2(n22307), .op(n17621) );
  and2_1 U19380 ( .ip1(n19236), .ip2(n17621), .op(n17622) );
  nor2_1 U19381 ( .ip1(n17623), .ip2(n17622), .op(n17624) );
  or2_1 U19382 ( .ip1(n22308), .ip2(n17624), .op(n17627) );
  or2_1 U19383 ( .ip1(n17625), .ip2(n17624), .op(n17626) );
  nand2_1 U19384 ( .ip1(n17627), .ip2(n17626), .op(\pipeline/csr/N1931 ) );
  inv_1 U19385 ( .ip(n17628), .op(n17629) );
  nand2_1 U19386 ( .ip1(n17630), .ip2(n17629), .op(n17651) );
  inv_1 U19387 ( .ip(n17651), .op(n17631) );
  and2_1 U19388 ( .ip1(n17632), .ip2(n17631), .op(n17633) );
  nor2_1 U19389 ( .ip1(n21089), .ip2(n17633), .op(n17634) );
  or2_1 U19390 ( .ip1(n17634), .ip2(n21120), .op(n22284) );
  inv_1 U19391 ( .ip(n22284), .op(n22276) );
  inv_1 U19392 ( .ip(\pipeline/csr/time_full [61]), .op(n18953) );
  inv_1 U19393 ( .ip(\pipeline/csr/time_full [59]), .op(n17650) );
  inv_1 U19394 ( .ip(\pipeline/csr/time_full [57]), .op(n18823) );
  inv_1 U19395 ( .ip(\pipeline/csr/time_full [55]), .op(n22278) );
  inv_1 U19396 ( .ip(\pipeline/csr/time_full [51]), .op(n18584) );
  inv_1 U19397 ( .ip(\pipeline/csr/time_full [49]), .op(n19973) );
  inv_1 U19398 ( .ip(\pipeline/csr/time_full [47]), .op(n19450) );
  inv_1 U19399 ( .ip(\pipeline/csr/time_full [45]), .op(n20252) );
  inv_1 U19400 ( .ip(\pipeline/csr/time_full [43]), .op(n20174) );
  inv_1 U19401 ( .ip(\pipeline/csr/time_full [41]), .op(n18436) );
  inv_1 U19402 ( .ip(\pipeline/csr/time_full [39]), .op(n19561) );
  inv_1 U19403 ( .ip(\pipeline/csr/time_full [35]), .op(n22271) );
  inv_1 U19404 ( .ip(\pipeline/csr/time_full [33]), .op(n22264) );
  inv_1 U19405 ( .ip(\pipeline/csr/time_full [31]), .op(n17648) );
  inv_1 U19406 ( .ip(\pipeline/csr/time_full [29]), .op(n17647) );
  inv_1 U19407 ( .ip(\pipeline/csr/time_full [27]), .op(n17646) );
  inv_1 U19408 ( .ip(\pipeline/csr/time_full [25]), .op(n17645) );
  inv_1 U19409 ( .ip(\pipeline/csr/time_full [23]), .op(n17644) );
  inv_1 U19410 ( .ip(\pipeline/csr/time_full [19]), .op(n17642) );
  inv_1 U19411 ( .ip(\pipeline/csr/time_full [17]), .op(n17641) );
  inv_1 U19412 ( .ip(\pipeline/csr/time_full [15]), .op(n17640) );
  inv_1 U19413 ( .ip(\pipeline/csr/time_full [13]), .op(n17639) );
  inv_1 U19414 ( .ip(\pipeline/csr/time_full [11]), .op(n20184) );
  inv_1 U19415 ( .ip(\pipeline/csr/time_full [9]), .op(n17638) );
  inv_1 U19416 ( .ip(\pipeline/csr/time_full [7]), .op(n17637) );
  inv_1 U19417 ( .ip(\pipeline/csr/time_full [5]), .op(n17636) );
  inv_1 U19418 ( .ip(\pipeline/csr/time_full [3]), .op(n17635) );
  nand3_1 U19419 ( .ip1(\pipeline/csr/time_full [2]), .ip2(
        \pipeline/csr/time_full [1]), .ip3(\pipeline/csr/time_full [0]), .op(
        n21175) );
  nor2_1 U19420 ( .ip1(n17635), .ip2(n21175), .op(n21180) );
  nand2_1 U19421 ( .ip1(\pipeline/csr/time_full [4]), .ip2(n21180), .op(n21055) );
  nor2_1 U19422 ( .ip1(n17636), .ip2(n21055), .op(n21058) );
  nand2_1 U19423 ( .ip1(\pipeline/csr/time_full [6]), .ip2(n21058), .op(n20344) );
  nor2_1 U19424 ( .ip1(n17637), .ip2(n20344), .op(n19702) );
  nand2_1 U19425 ( .ip1(\pipeline/csr/time_full [8]), .ip2(n19702), .op(n18428) );
  nor2_1 U19426 ( .ip1(n17638), .ip2(n18428), .op(n19784) );
  nand2_1 U19427 ( .ip1(\pipeline/csr/time_full [10]), .ip2(n19784), .op(
        n20183) );
  nor2_1 U19428 ( .ip1(n20184), .ip2(n20183), .op(n20752) );
  nand2_1 U19429 ( .ip1(\pipeline/csr/time_full [12]), .ip2(n20752), .op(
        n20754) );
  nor2_1 U19430 ( .ip1(n17639), .ip2(n20754), .op(n20246) );
  nand2_1 U19431 ( .ip1(\pipeline/csr/time_full [14]), .ip2(n20246), .op(
        n19851) );
  nor2_1 U19432 ( .ip1(n17640), .ip2(n19851), .op(n19909) );
  nand2_1 U19433 ( .ip1(\pipeline/csr/time_full [16]), .ip2(n19909), .op(
        n19977) );
  nor2_1 U19434 ( .ip1(n17641), .ip2(n19977), .op(n19980) );
  nand2_1 U19435 ( .ip1(\pipeline/csr/time_full [18]), .ip2(n19980), .op(
        n18588) );
  nor2_1 U19436 ( .ip1(n17642), .ip2(n18588), .op(n19512) );
  nand2_1 U19437 ( .ip1(\pipeline/csr/time_full [20]), .ip2(n19512), .op(
        n18655) );
  nor2_1 U19438 ( .ip1(n17643), .ip2(n18655), .op(n20063) );
  nand2_1 U19439 ( .ip1(\pipeline/csr/time_full [22]), .ip2(n20063), .op(
        n20115) );
  nor2_1 U19440 ( .ip1(n17644), .ip2(n20115), .op(n20118) );
  nand2_1 U19441 ( .ip1(\pipeline/csr/time_full [24]), .ip2(n20118), .op(
        n18757) );
  nor2_1 U19442 ( .ip1(n17645), .ip2(n18757), .op(n19097) );
  nand2_1 U19443 ( .ip1(\pipeline/csr/time_full [26]), .ip2(n19097), .op(
        n19216) );
  nor2_1 U19444 ( .ip1(n17646), .ip2(n19216), .op(n19254) );
  nand2_1 U19445 ( .ip1(\pipeline/csr/time_full [28]), .ip2(n19254), .op(
        n19256) );
  nor2_1 U19446 ( .ip1(n17647), .ip2(n19256), .op(n22251) );
  nand2_1 U19447 ( .ip1(\pipeline/csr/time_full [30]), .ip2(n22251), .op(
        n20924) );
  nor2_1 U19448 ( .ip1(n17648), .ip2(n20924), .op(n20927) );
  nand2_1 U19449 ( .ip1(\pipeline/csr/time_full [32]), .ip2(n20927), .op(
        n22263) );
  nor2_1 U19450 ( .ip1(n22264), .ip2(n22263), .op(n22262) );
  nand2_1 U19451 ( .ip1(\pipeline/csr/time_full [34]), .ip2(n22262), .op(
        n22270) );
  nor2_1 U19452 ( .ip1(n22271), .ip2(n22270), .op(n22269) );
  nand2_1 U19453 ( .ip1(\pipeline/csr/time_full [36]), .ip2(n22269), .op(
        n21052) );
  nor2_1 U19454 ( .ip1(n21051), .ip2(n21052), .op(n21050) );
  nand2_1 U19455 ( .ip1(\pipeline/csr/time_full [38]), .ip2(n21050), .op(
        n20330) );
  nor2_1 U19456 ( .ip1(n19561), .ip2(n20330), .op(n19695) );
  nand2_1 U19457 ( .ip1(\pipeline/csr/time_full [40]), .ip2(n19695), .op(
        n19697) );
  nor2_1 U19458 ( .ip1(n18436), .ip2(n19697), .op(n19780) );
  nand2_1 U19459 ( .ip1(\pipeline/csr/time_full [42]), .ip2(n19780), .op(
        n20175) );
  nor2_1 U19460 ( .ip1(n20174), .ip2(n20175), .op(n20747) );
  nand2_1 U19461 ( .ip1(\pipeline/csr/time_full [44]), .ip2(n20747), .op(
        n20253) );
  nor2_1 U19462 ( .ip1(n20252), .ip2(n20253), .op(n20251) );
  nand2_1 U19463 ( .ip1(\pipeline/csr/time_full [46]), .ip2(n20251), .op(
        n19847) );
  nor2_1 U19464 ( .ip1(n19450), .ip2(n19847), .op(n19449) );
  nand2_1 U19465 ( .ip1(\pipeline/csr/time_full [48]), .ip2(n19449), .op(
        n19974) );
  nor2_1 U19466 ( .ip1(n19973), .ip2(n19974), .op(n19972) );
  nand2_1 U19467 ( .ip1(\pipeline/csr/time_full [50]), .ip2(n19972), .op(
        n18585) );
  nor2_1 U19468 ( .ip1(n18584), .ip2(n18585), .op(n19508) );
  nand2_1 U19469 ( .ip1(\pipeline/csr/time_full [52]), .ip2(n19508), .op(
        n18651) );
  nor2_1 U19470 ( .ip1(n17649), .ip2(n18651), .op(n20059) );
  nand2_1 U19471 ( .ip1(\pipeline/csr/time_full [54]), .ip2(n20059), .op(
        n22277) );
  nor2_1 U19472 ( .ip1(n22278), .ip2(n22277), .op(n22275) );
  nand2_1 U19473 ( .ip1(\pipeline/csr/time_full [56]), .ip2(n22275), .op(
        n18824) );
  nor2_1 U19474 ( .ip1(n18823), .ip2(n18824), .op(n19093) );
  nand2_1 U19475 ( .ip1(\pipeline/csr/time_full [58]), .ip2(n19093), .op(
        n19239) );
  nor2_1 U19476 ( .ip1(n17650), .ip2(n19239), .op(n22283) );
  nand2_1 U19477 ( .ip1(\pipeline/csr/time_full [60]), .ip2(n22283), .op(
        n22286) );
  nor2_1 U19478 ( .ip1(n18953), .ip2(n22286), .op(n18952) );
  nand2_1 U19479 ( .ip1(\pipeline/csr/time_full [62]), .ip2(n18952), .op(
        n18881) );
  nor2_1 U19480 ( .ip1(\pipeline/csr/time_full [63]), .ip2(n18881), .op(n17653) );
  nor2_1 U19481 ( .ip1(n21089), .ip2(n17651), .op(n18435) );
  nand2_1 U19482 ( .ip1(n18435), .ip2(n20959), .op(n17655) );
  nor2_1 U19483 ( .ip1(n21210), .ip2(n17655), .op(n17652) );
  not_ab_or_c_or_d U19484 ( .ip1(\pipeline/csr/time_full [63]), .ip2(n18881), 
        .ip3(n17653), .ip4(n17652), .op(n17654) );
  or2_1 U19485 ( .ip1(n22276), .ip2(n17654), .op(n17657) );
  or2_1 U19486 ( .ip1(n17655), .ip2(n17654), .op(n17656) );
  nand2_1 U19487 ( .ip1(n17657), .ip2(n17656), .op(\pipeline/csr/N2000 ) );
  nand2_1 U19488 ( .ip1(n18435), .ip2(n19951), .op(n17662) );
  nor2_1 U19489 ( .ip1(n21210), .ip2(n17662), .op(n17660) );
  or2_1 U19490 ( .ip1(\pipeline/csr/time_full [48]), .ip2(n19449), .op(n17658)
         );
  and2_1 U19491 ( .ip1(n19974), .ip2(n17658), .op(n17659) );
  nor2_1 U19492 ( .ip1(n17660), .ip2(n17659), .op(n17661) );
  or2_1 U19493 ( .ip1(n22276), .ip2(n17661), .op(n17664) );
  or2_1 U19494 ( .ip1(n17662), .ip2(n17661), .op(n17663) );
  nand2_1 U19495 ( .ip1(n17664), .ip2(n17663), .op(\pipeline/csr/N1985 ) );
  inv_1 U19496 ( .ip(n17665), .op(n17667) );
  inv_1 U19497 ( .ip(n17666), .op(n21528) );
  nor2_1 U19498 ( .ip1(n17667), .ip2(n21528), .op(n17668) );
  nand2_1 U19499 ( .ip1(n21531), .ip2(n17668), .op(n17670) );
  and2_1 U19500 ( .ip1(n17670), .ip2(n17669), .op(n17806) );
  nor2_1 U19501 ( .ip1(imem_hready), .ip2(n10364), .op(n17671) );
  nand2_1 U19502 ( .ip1(n17806), .ip2(n17671), .op(n17672) );
  nand2_1 U19503 ( .ip1(n17672), .ip2(n17816), .op(n17790) );
  or2_1 U19504 ( .ip1(n21089), .ip2(n17790), .op(n19766) );
  inv_1 U19505 ( .ip(n19766), .op(n21995) );
  nand2_1 U19506 ( .ip1(imem_hready), .ip2(imem_badmem_e), .op(n17803) );
  and3_1 U19507 ( .ip1(n17674), .ip2(n17673), .ip3(n17803), .op(n17675) );
  and2_1 U19508 ( .ip1(n17806), .ip2(n17675), .op(n17676) );
  and2_1 U19509 ( .ip1(n21995), .ip2(n17676), .op(n21988) );
  inv_1 U19510 ( .ip(n21988), .op(n17680) );
  or2_1 U19511 ( .ip1(htif_reset), .ip2(n17816), .op(n17677) );
  nand2_1 U19512 ( .ip1(n17680), .ip2(n17677), .op(n17691) );
  inv_1 U19513 ( .ip(n17677), .op(n22049) );
  nand2_1 U19514 ( .ip1(\pipeline/inst_DX [0]), .ip2(n22049), .op(n17679) );
  nand2_1 U19515 ( .ip1(n21988), .ip2(imem_rdata[0]), .op(n17678) );
  nand3_1 U19516 ( .ip1(n17691), .ip2(n17679), .ip3(n17678), .op(n8503) );
  inv_1 U19517 ( .ip(n17680), .op(n22048) );
  nand2_1 U19518 ( .ip1(n22048), .ip2(imem_rdata[1]), .op(n17682) );
  nand2_1 U19519 ( .ip1(\pipeline/inst_DX [1]), .ip2(n22049), .op(n17681) );
  nand3_1 U19520 ( .ip1(n17691), .ip2(n17682), .ip3(n17681), .op(n8502) );
  nand2_1 U19521 ( .ip1(n22048), .ip2(imem_rdata[13]), .op(n17684) );
  nand2_1 U19522 ( .ip1(dmem_hsize[1]), .ip2(n22049), .op(n17683) );
  nand2_1 U19523 ( .ip1(n17684), .ip2(n17683), .op(n8523) );
  nand2_1 U19524 ( .ip1(n22048), .ip2(imem_rdata[14]), .op(n17686) );
  nand2_1 U19525 ( .ip1(\pipeline/dmem_type[2] ), .ip2(n22049), .op(n17685) );
  nand2_1 U19526 ( .ip1(n17686), .ip2(n17685), .op(n8522) );
  nand2_1 U19527 ( .ip1(n21988), .ip2(imem_rdata[12]), .op(n17688) );
  nand2_1 U19528 ( .ip1(dmem_hsize[0]), .ip2(n22049), .op(n17687) );
  nand2_1 U19529 ( .ip1(n17688), .ip2(n17687), .op(n8524) );
  nand2_1 U19530 ( .ip1(n21988), .ip2(imem_rdata[4]), .op(n17690) );
  nand2_1 U19531 ( .ip1(\pipeline/inst_DX [4]), .ip2(n22049), .op(n17689) );
  nand3_1 U19532 ( .ip1(n17691), .ip2(n17690), .ip3(n17689), .op(n8501) );
  nand2_1 U19533 ( .ip1(n22048), .ip2(imem_rdata[6]), .op(n17693) );
  nand2_1 U19534 ( .ip1(\pipeline/inst_DX [6]), .ip2(n22049), .op(n17692) );
  nand2_1 U19535 ( .ip1(n17693), .ip2(n17692), .op(n8530) );
  nand2_1 U19536 ( .ip1(n21988), .ip2(imem_rdata[5]), .op(n17695) );
  nand2_1 U19537 ( .ip1(\pipeline/inst_DX [5]), .ip2(n22049), .op(n17694) );
  nand2_1 U19538 ( .ip1(n17695), .ip2(n17694), .op(n8531) );
  nand2_1 U19539 ( .ip1(n22048), .ip2(imem_rdata[2]), .op(n17697) );
  nand2_1 U19540 ( .ip1(\pipeline/inst_DX [2]), .ip2(n22049), .op(n17696) );
  nand2_1 U19541 ( .ip1(n17697), .ip2(n17696), .op(n8533) );
  nand2_1 U19542 ( .ip1(n22048), .ip2(imem_rdata[3]), .op(n17699) );
  nand2_1 U19543 ( .ip1(\pipeline/inst_DX [3]), .ip2(n22049), .op(n17698) );
  nand2_1 U19544 ( .ip1(n17699), .ip2(n17698), .op(n8532) );
  nand2_1 U19545 ( .ip1(n22048), .ip2(imem_rdata[15]), .op(n17701) );
  nand2_1 U19546 ( .ip1(\pipeline/inst_DX [15]), .ip2(n22049), .op(n17700) );
  nand2_1 U19547 ( .ip1(n17701), .ip2(n17700), .op(n8520) );
  nand2_1 U19548 ( .ip1(n22048), .ip2(imem_rdata[16]), .op(n17703) );
  nand2_1 U19549 ( .ip1(\pipeline/inst_DX [16]), .ip2(n22049), .op(n17702) );
  nand2_1 U19550 ( .ip1(n17703), .ip2(n17702), .op(n8519) );
  nand2_1 U19551 ( .ip1(n21988), .ip2(imem_rdata[18]), .op(n17705) );
  nand2_1 U19552 ( .ip1(\pipeline/inst_DX [18]), .ip2(n22049), .op(n17704) );
  nand2_1 U19553 ( .ip1(n17705), .ip2(n17704), .op(n8517) );
  nand2_1 U19554 ( .ip1(n22048), .ip2(imem_rdata[19]), .op(n17707) );
  nand2_1 U19555 ( .ip1(\pipeline/inst_DX [19]), .ip2(n22049), .op(n17706) );
  nand2_1 U19556 ( .ip1(n17707), .ip2(n17706), .op(n8516) );
  nand2_1 U19557 ( .ip1(n21988), .ip2(imem_rdata[17]), .op(n17709) );
  nand2_1 U19558 ( .ip1(\pipeline/inst_DX [17]), .ip2(n22049), .op(n17708) );
  nand2_1 U19559 ( .ip1(n17709), .ip2(n17708), .op(n8518) );
  nand2_1 U19560 ( .ip1(n21988), .ip2(imem_rdata[11]), .op(n17711) );
  nand2_1 U19561 ( .ip1(\pipeline/inst_DX [11]), .ip2(n22049), .op(n17710) );
  nand2_1 U19562 ( .ip1(n17711), .ip2(n17710), .op(n8525) );
  nand2_1 U19563 ( .ip1(n22048), .ip2(imem_rdata[10]), .op(n17713) );
  nand2_1 U19564 ( .ip1(\pipeline/inst_DX [10]), .ip2(n22049), .op(n17712) );
  nand2_1 U19565 ( .ip1(n17713), .ip2(n17712), .op(n8526) );
  nand2_1 U19566 ( .ip1(n22048), .ip2(imem_rdata[9]), .op(n17715) );
  nand2_1 U19567 ( .ip1(\pipeline/inst_DX [9]), .ip2(n22049), .op(n17714) );
  nand2_1 U19568 ( .ip1(n17715), .ip2(n17714), .op(n8527) );
  nand2_1 U19569 ( .ip1(n22048), .ip2(imem_rdata[8]), .op(n17717) );
  nand2_1 U19570 ( .ip1(\pipeline/inst_DX [8]), .ip2(n22049), .op(n17716) );
  nand2_1 U19571 ( .ip1(n17717), .ip2(n17716), .op(n8528) );
  nand2_1 U19572 ( .ip1(n22048), .ip2(imem_rdata[7]), .op(n17719) );
  nand2_1 U19573 ( .ip1(\pipeline/inst_DX [7]), .ip2(n22049), .op(n17718) );
  nand2_1 U19574 ( .ip1(n17719), .ip2(n17718), .op(n8529) );
  nand2_1 U19575 ( .ip1(n21988), .ip2(imem_rdata[26]), .op(n17721) );
  nand2_1 U19576 ( .ip1(\pipeline/inst_DX [26]), .ip2(n22049), .op(n17720) );
  nand2_1 U19577 ( .ip1(n17721), .ip2(n17720), .op(n8509) );
  nand2_1 U19578 ( .ip1(n21988), .ip2(imem_rdata[22]), .op(n17723) );
  nand2_1 U19579 ( .ip1(\pipeline/inst_DX [22]), .ip2(n22049), .op(n17722) );
  nand2_1 U19580 ( .ip1(n17723), .ip2(n17722), .op(n8513) );
  nand2_1 U19581 ( .ip1(n22048), .ip2(imem_rdata[24]), .op(n17725) );
  nand2_1 U19582 ( .ip1(\pipeline/inst_DX [24]), .ip2(n22049), .op(n17724) );
  nand2_1 U19583 ( .ip1(n17725), .ip2(n17724), .op(n8511) );
  nand2_1 U19584 ( .ip1(n22048), .ip2(imem_rdata[23]), .op(n17727) );
  nand2_1 U19585 ( .ip1(\pipeline/inst_DX [23]), .ip2(n22049), .op(n17726) );
  nand2_1 U19586 ( .ip1(n17727), .ip2(n17726), .op(n8512) );
  nand2_1 U19587 ( .ip1(n22048), .ip2(imem_rdata[29]), .op(n17729) );
  nand2_1 U19588 ( .ip1(\pipeline/inst_DX [29]), .ip2(n22049), .op(n17728) );
  nand2_1 U19589 ( .ip1(n17729), .ip2(n17728), .op(n8506) );
  nand2_1 U19590 ( .ip1(n22048), .ip2(imem_rdata[31]), .op(n17731) );
  nand2_1 U19591 ( .ip1(\pipeline/imm[31] ), .ip2(n22049), .op(n17730) );
  nand2_1 U19592 ( .ip1(n17731), .ip2(n17730), .op(n8504) );
  nand2_1 U19593 ( .ip1(n21988), .ip2(imem_rdata[27]), .op(n17733) );
  nand2_1 U19594 ( .ip1(\pipeline/inst_DX [27]), .ip2(n22049), .op(n17732) );
  nand2_1 U19595 ( .ip1(n17733), .ip2(n17732), .op(n8508) );
  nand2_1 U19596 ( .ip1(n21988), .ip2(imem_rdata[21]), .op(n17735) );
  nand2_1 U19597 ( .ip1(\pipeline/inst_DX [21]), .ip2(n22049), .op(n17734) );
  nand2_1 U19598 ( .ip1(n17735), .ip2(n17734), .op(n8514) );
  nand2_1 U19599 ( .ip1(n22048), .ip2(imem_rdata[20]), .op(n17737) );
  nand2_1 U19600 ( .ip1(\pipeline/inst_DX [20]), .ip2(n22049), .op(n17736) );
  nand2_1 U19601 ( .ip1(n17737), .ip2(n17736), .op(n8515) );
  nand2_1 U19602 ( .ip1(n22048), .ip2(imem_rdata[28]), .op(n17739) );
  nand2_1 U19603 ( .ip1(\pipeline/inst_DX [28]), .ip2(n22049), .op(n17738) );
  nand2_1 U19604 ( .ip1(n17739), .ip2(n17738), .op(n8507) );
  nor2_1 U19605 ( .ip1(n17740), .ip2(n17819), .op(dmem_htrans[1]) );
  inv_1 U19606 ( .ip(dmem_htrans[1]), .op(n17887) );
  nor2_1 U19607 ( .ip1(n17784), .ip2(n17887), .op(dmem_hwrite) );
  buf_1 U19608 ( .ip(n21582), .op(n19505) );
  nand2_1 U19609 ( .ip1(n22067), .ip2(dmem_hwrite), .op(n17743) );
  nor2_1 U19610 ( .ip1(htif_reset), .ip2(n17741), .op(n22043) );
  nand2_1 U19611 ( .ip1(\pipeline/ctrl/store_in_WB ), .ip2(n22043), .op(n17742) );
  nand2_1 U19612 ( .ip1(n17743), .ip2(n17742), .op(n8498) );
  inv_1 U19613 ( .ip(imem_hready), .op(n17746) );
  inv_1 U19614 ( .ip(n17806), .op(n17745) );
  ab_or_c_or_d U19615 ( .ip1(n17746), .ip2(n17745), .ip3(n17744), .ip4(n21089), 
        .op(\pipeline/ctrl/N66 ) );
  nand2_1 U19616 ( .ip1(n21440), .ip2(n17747), .op(n17762) );
  nor3_1 U19617 ( .ip1(n21493), .ip2(\pipeline/md/counter [2]), .ip3(n18213), 
        .op(n17758) );
  ab_or_c_or_d U19618 ( .ip1(\pipeline/md/counter [2]), .ip2(n17762), .ip3(
        n22042), .ip4(n17758), .op(n8536) );
  nand2_1 U19619 ( .ip1(n14765), .ip2(n17751), .op(n17748) );
  nor2_1 U19620 ( .ip1(\pipeline/md/counter [4]), .ip2(n17748), .op(n17749) );
  ab_or_c_or_d U19621 ( .ip1(\pipeline/md/counter [4]), .ip2(n17748), .ip3(
        n22042), .ip4(n17749), .op(n8534) );
  nor2_1 U19622 ( .ip1(n20552), .ip2(n17749), .op(n17750) );
  nor2_1 U19623 ( .ip1(htif_reset), .ip2(n17750), .op(\pipeline/md/N162 ) );
  inv_1 U19624 ( .ip(n17751), .op(n21516) );
  nor2_1 U19625 ( .ip1(\pipeline/md/counter [4]), .ip2(n21516), .op(n17752) );
  nor2_1 U19626 ( .ip1(n17752), .ip2(n22665), .op(n17753) );
  nor2_1 U19627 ( .ip1(n20552), .ip2(n17753), .op(n17754) );
  nand2_1 U19628 ( .ip1(n21683), .ip2(n17754), .op(n17755) );
  xor2_1 U19629 ( .ip1(\pipeline/md/counter [0]), .ip2(n22665), .op(n17757) );
  nand2_1 U19630 ( .ip1(n21683), .ip2(n17757), .op(n8538) );
  nor2_1 U19631 ( .ip1(\pipeline/md/counter [3]), .ip2(n17758), .op(n17759) );
  nor2_1 U19632 ( .ip1(n17760), .ip2(n17759), .op(n17761) );
  ab_or_c_or_d U19633 ( .ip1(\pipeline/md/counter [3]), .ip2(n17762), .ip3(
        n22042), .ip4(n17761), .op(n8535) );
  nand3_1 U19634 ( .ip1(dmem_hsize[1]), .ip2(\pipeline/dmem_type[2] ), .ip3(
        n22042), .op(n17769) );
  nand2_1 U19635 ( .ip1(\pipeline/md/op [1]), .ip2(n21683), .op(n17763) );
  nand2_1 U19636 ( .ip1(n17769), .ip2(n17763), .op(n10061) );
  nor2_1 U19637 ( .ip1(dmem_hsize[1]), .ip2(n17765), .op(n17764) );
  mux2_1 U19638 ( .ip1(\pipeline/md/op [0]), .ip2(n17764), .s(n22042), .op(
        n10062) );
  inv_1 U19639 ( .ip(n21582), .op(n19498) );
  mux2_1 U19640 ( .ip1(\pipeline/dmem_type_WB [1]), .ip2(dmem_hsize[1]), .s(
        n17429), .op(n8774) );
  mux2_1 U19641 ( .ip1(\pipeline/dmem_type_WB [2]), .ip2(
        \pipeline/dmem_type[2] ), .s(n17777), .op(n8773) );
  nand3_1 U19642 ( .ip1(n22042), .ip2(n17765), .ip3(n22090), .op(n17767) );
  nand2_1 U19643 ( .ip1(\pipeline/md/out_sel [0]), .ip2(n21683), .op(n17766)
         );
  nand2_1 U19644 ( .ip1(n17767), .ip2(n17766), .op(n10064) );
  nand2_1 U19645 ( .ip1(\pipeline/md/out_sel [1]), .ip2(n21683), .op(n17768)
         );
  nand2_1 U19646 ( .ip1(n17769), .ip2(n17768), .op(n10063) );
  inv_1 U19647 ( .ip(\pipeline/md/op [1]), .op(n17770) );
  nor2_1 U19648 ( .ip1(\pipeline/md/op [0]), .ip2(n17770), .op(n17771) );
  nor3_1 U19649 ( .ip1(n21624), .ip2(n17771), .ip3(n21406), .op(n17776) );
  inv_1 U19650 ( .ip(n17771), .op(n17772) );
  nor2_1 U19651 ( .ip1(n21683), .ip2(n17772), .op(n17773) );
  nor2_1 U19652 ( .ip1(n21400), .ip2(n17773), .op(n17774) );
  nor2_1 U19653 ( .ip1(n17774), .ip2(n20483), .op(n17775) );
  ab_or_c_or_d U19654 ( .ip1(\pipeline/md/negate_output ), .ip2(n21683), .ip3(
        n17776), .ip4(n17775), .op(n8904) );
  nand2_1 U19655 ( .ip1(\pipeline/ctrl/wfi_unkilled_WB ), .ip2(n22043), .op(
        n17781) );
  inv_1 U19656 ( .ip(n21582), .op(n17777) );
  nand4_1 U19657 ( .ip1(n17779), .ip2(n17778), .ip3(n17891), .ip4(n20389), 
        .op(n17780) );
  nand2_1 U19658 ( .ip1(n17781), .ip2(n17780), .op(n8494) );
  nand2_1 U19659 ( .ip1(n17788), .ip2(n17782), .op(n17783) );
  mux2_1 U19660 ( .ip1(\pipeline/wb_src_sel_WB [1]), .ip2(n17783), .s(n17777), 
        .op(n10065) );
  nand3_1 U19661 ( .ip1(n17786), .ip2(n17785), .ip3(n17784), .op(n17787) );
  nand2_1 U19662 ( .ip1(n17788), .ip2(n17787), .op(n17789) );
  mux2_1 U19663 ( .ip1(\pipeline/wb_src_sel_WB [0]), .ip2(n17789), .s(n22067), 
        .op(n10066) );
  nand2_1 U19664 ( .ip1(n21995), .ip2(imem_haddr[2]), .op(n17792) );
  nand2_1 U19665 ( .ip1(n17790), .ip2(n20966), .op(n19765) );
  inv_1 U19666 ( .ip(n19765), .op(n21996) );
  nand2_1 U19667 ( .ip1(\pipeline/PC_IF [2]), .ip2(n21996), .op(n17791) );
  nand2_1 U19668 ( .ip1(n17792), .ip2(n17791), .op(n8486) );
  nand2_1 U19669 ( .ip1(\pipeline/PC_IF [2]), .ip2(n21988), .op(n17794) );
  or2_1 U19670 ( .ip1(htif_reset), .ip2(n21988), .op(n17817) );
  inv_1 U19671 ( .ip(n17817), .op(n21999) );
  nand2_1 U19672 ( .ip1(\pipeline/PC_DX [2]), .ip2(n21999), .op(n17793) );
  nand2_1 U19673 ( .ip1(n17794), .ip2(n17793), .op(n8485) );
  mux2_1 U19674 ( .ip1(\pipeline/PC_WB [2]), .ip2(\pipeline/PC_DX [2]), .s(
        n19498), .op(n8901) );
  nand2_1 U19675 ( .ip1(n22351), .ip2(n21043), .op(n17798) );
  inv_1 U19676 ( .ip(n21171), .op(n21046) );
  xor2_1 U19677 ( .ip1(\pipeline/PC_WB [2]), .ip2(n20972), .op(n17795) );
  nand2_1 U19678 ( .ip1(n21046), .ip2(n17795), .op(n17797) );
  nand2_1 U19679 ( .ip1(n21174), .ip2(\pipeline/epc [2]), .op(n17796) );
  nand3_1 U19680 ( .ip1(n17798), .ip2(n17797), .ip3(n17796), .op(n8869) );
  nor2_1 U19681 ( .ip1(n22351), .ip2(n21029), .op(n17802) );
  nor2_1 U19682 ( .ip1(htif_reset), .ip2(n21029), .op(n21032) );
  inv_1 U19683 ( .ip(\pipeline/csr/mtvec [2]), .op(n17799) );
  nor2_1 U19684 ( .ip1(htif_reset), .ip2(n17799), .op(n17800) );
  nor2_1 U19685 ( .ip1(n21032), .ip2(n17800), .op(n17801) );
  nor2_1 U19686 ( .ip1(n17802), .ip2(n17801), .op(n9990) );
  nand2_1 U19687 ( .ip1(\pipeline/ctrl/had_ex_DX ), .ip2(n22049), .op(n17808)
         );
  nor4_1 U19688 ( .ip1(n21089), .ip2(\pipeline/ctrl/replay_IF ), .ip3(n17804), 
        .ip4(n17803), .op(n17805) );
  nand2_1 U19689 ( .ip1(n17806), .ip2(n17805), .op(n17807) );
  nand2_1 U19690 ( .ip1(n17808), .ip2(n17807), .op(n8500) );
  nand2_1 U19691 ( .ip1(n21032), .ip2(n22145), .op(n17811) );
  inv_1 U19692 ( .ip(n21029), .op(n17809) );
  nor2_1 U19693 ( .ip1(htif_reset), .ip2(n17809), .op(n20705) );
  nand2_1 U19694 ( .ip1(\pipeline/csr/mtvec [5]), .ip2(n20705), .op(n17810) );
  nand2_1 U19695 ( .ip1(n17811), .ip2(n17810), .op(n9987) );
  nand2_1 U19696 ( .ip1(n17812), .ip2(n20965), .op(n22371) );
  inv_1 U19697 ( .ip(n22371), .op(n17813) );
  nor2_1 U19698 ( .ip1(htif_reset), .ip2(n17813), .op(n22363) );
  nand2_1 U19699 ( .ip1(\pipeline/csr/mtimecmp [5]), .ip2(n22363), .op(n17815)
         );
  nor2_1 U19700 ( .ip1(htif_reset), .ip2(n22371), .op(n22365) );
  nand2_1 U19701 ( .ip1(n22365), .ip2(n22145), .op(n17814) );
  nand2_1 U19702 ( .ip1(n17815), .ip2(n17814), .op(n10017) );
  nor2_1 U19703 ( .ip1(n17816), .ip2(\pipeline/ctrl/prev_killed_DX ), .op(
        n17818) );
  nor2_1 U19704 ( .ip1(n17818), .ip2(n17817), .op(n8492) );
  nand2_1 U19705 ( .ip1(\pipeline/ctrl/prev_killed_WB ), .ip2(n22043), .op(
        n17822) );
  or2_1 U19706 ( .ip1(\pipeline/ctrl/prev_killed_DX ), .ip2(n17819), .op(
        n17820) );
  nand2_1 U19707 ( .ip1(n22067), .ip2(n17820), .op(n17821) );
  nand2_1 U19708 ( .ip1(n17822), .ip2(n17821), .op(n8491) );
  inv_1 U19709 ( .ip(n21001), .op(n21019) );
  inv_1 U19710 ( .ip(n21016), .op(n20990) );
  nor2_1 U19711 ( .ip1(n17824), .ip2(n20990), .op(n17827) );
  mux2_1 U19712 ( .ip1(n17824), .ip2(\pipeline/csr/instret_full [5]), .s(
        n17823), .op(n17825) );
  nor2_1 U19713 ( .ip1(n21005), .ip2(n17825), .op(n17826) );
  ab_or_c_or_d U19714 ( .ip1(n21019), .ip2(n22145), .ip3(n17827), .ip4(n17826), 
        .op(n10133) );
  nand2_1 U19715 ( .ip1(n17828), .ip2(n20965), .op(n17830) );
  inv_1 U19716 ( .ip(n17830), .op(n17829) );
  nor2_1 U19717 ( .ip1(htif_reset), .ip2(n17829), .op(n22013) );
  nand2_1 U19718 ( .ip1(\pipeline/csr/mscratch [5]), .ip2(n22013), .op(n17832)
         );
  nor2_1 U19719 ( .ip1(htif_reset), .ip2(n17830), .op(n22014) );
  nand2_1 U19720 ( .ip1(n22014), .ip2(n22145), .op(n17831) );
  nand2_1 U19721 ( .ip1(n17832), .ip2(n17831), .op(n9923) );
  inv_1 U19722 ( .ip(n20965), .op(n19601) );
  nor2_1 U19723 ( .ip1(n19601), .ip2(n17833), .op(n17834) );
  nor2_1 U19724 ( .ip1(htif_reset), .ip2(n17834), .op(n22372) );
  nand2_1 U19725 ( .ip1(\pipeline/csr/from_host [5]), .ip2(n22372), .op(n17837) );
  inv_1 U19726 ( .ip(n17834), .op(n17835) );
  nor2_1 U19727 ( .ip1(htif_reset), .ip2(n17835), .op(n22373) );
  nand2_1 U19728 ( .ip1(n22373), .ip2(n22145), .op(n17836) );
  nand2_1 U19729 ( .ip1(n17837), .ip2(n17836), .op(n9955) );
  nand3_1 U19730 ( .ip1(htif_pcr_req_addr[9]), .ip2(htif_pcr_req_addr[8]), 
        .ip3(htif_pcr_req_addr[10]), .op(n17838) );
  nor2_1 U19731 ( .ip1(htif_pcr_req_addr[11]), .ip2(n17838), .op(n17841) );
  nor3_1 U19732 ( .ip1(htif_pcr_req_addr[5]), .ip2(htif_pcr_req_addr[1]), 
        .ip3(htif_pcr_req_addr[3]), .op(n17840) );
  nor4_1 U19733 ( .ip1(htif_pcr_req_addr[4]), .ip2(htif_pcr_req_addr[2]), 
        .ip3(htif_pcr_req_addr[6]), .ip4(n22476), .op(n17839) );
  nand4_1 U19734 ( .ip1(n17841), .ip2(htif_pcr_req_addr[7]), .ip3(n17840), 
        .ip4(n17839), .op(n22381) );
  nor2_1 U19735 ( .ip1(htif_pcr_req_addr[0]), .ip2(n22381), .op(n22477) );
  inv_1 U19736 ( .ip(\pipeline/csr/system_wen ), .op(n17847) );
  nand2_1 U19737 ( .ip1(n22477), .ip2(n17847), .op(n17842) );
  nand2_1 U19738 ( .ip1(n20966), .ip2(n17842), .op(n17845) );
  nor2_1 U19739 ( .ip1(n19601), .ip2(n17843), .op(n17846) );
  inv_1 U19740 ( .ip(n17846), .op(n17844) );
  nor2_1 U19741 ( .ip1(n17845), .ip2(n17844), .op(n22378) );
  nand2_1 U19742 ( .ip1(n22378), .ip2(n22145), .op(n17849) );
  not_ab_or_c_or_d U19743 ( .ip1(n22477), .ip2(n17847), .ip3(n17846), .ip4(
        n21089), .op(n22376) );
  nand2_1 U19744 ( .ip1(\pipeline/csr/to_host [5]), .ip2(n22376), .op(n17848)
         );
  nand2_1 U19745 ( .ip1(n17849), .ip2(n17848), .op(n8767) );
  fulladder U19746 ( .a(\pipeline/md/a [3]), .b(n17851), .ci(n17850), .co(
        n14651), .s(n17852) );
  nand2_1 U19747 ( .ip1(n21944), .ip2(n17852), .op(n17859) );
  buf_1 U19748 ( .ip(n21947), .op(n21884) );
  nand2_1 U19749 ( .ip1(n21884), .ip2(\pipeline/md/a [3]), .op(n17858) );
  nand2_1 U19750 ( .ip1(n21624), .ip2(n17853), .op(n17854) );
  xor2_1 U19751 ( .ip1(n17855), .ip2(n17854), .op(n17856) );
  nand2_1 U19752 ( .ip1(n21649), .ip2(n17856), .op(n17857) );
  nand3_1 U19753 ( .ip1(n17859), .ip2(n17858), .ip3(n17857), .op(n8380) );
  nand2_1 U19754 ( .ip1(n17861), .ip2(n17860), .op(n17862) );
  nand2_1 U19755 ( .ip1(n14765), .ip2(n17862), .op(n17863) );
  nand2_1 U19756 ( .ip1(n22738), .ip2(n17863), .op(n17879) );
  nor3_1 U19757 ( .ip1(n17865), .ip2(n22755), .ip3(n17864), .op(n17878) );
  nand2_1 U19758 ( .ip1(\pipeline/md/negate_output ), .ip2(n17866), .op(n17868) );
  nor2_1 U19759 ( .ip1(n17869), .ip2(n17868), .op(n17867) );
  not_ab_or_c_or_d U19760 ( .ip1(n17869), .ip2(n17868), .ip3(n17867), .ip4(
        n21960), .op(n17876) );
  inv_1 U19761 ( .ip(\pipeline/md/result [35]), .op(n22519) );
  nor2_1 U19762 ( .ip1(n21967), .ip2(n22519), .op(n17870) );
  not_ab_or_c_or_d U19763 ( .ip1(n17872), .ip2(n17871), .ip3(n21972), .ip4(
        n17870), .op(n17875) );
  nor3_1 U19764 ( .ip1(n22519), .ip2(n17873), .ip3(n21505), .op(n17874) );
  nor3_1 U19765 ( .ip1(n17876), .ip2(n17875), .ip3(n17874), .op(n17877) );
  not_ab_or_c_or_d U19766 ( .ip1(\pipeline/md_resp_result [3]), .ip2(n17879), 
        .ip3(n17878), .ip4(n17877), .op(n17881) );
  nand2_1 U19767 ( .ip1(n20554), .ip2(n21271), .op(n17880) );
  nand2_1 U19768 ( .ip1(n17881), .ip2(n17880), .op(n8631) );
  mux2_1 U19769 ( .ip1(\pipeline/csr_rdata_WB [3]), .ip2(n17882), .s(n22067), 
        .op(n8803) );
  mux2_1 U19770 ( .ip1(\pipeline/reg_to_wr_WB [0]), .ip2(\pipeline/inst_DX [7]), .s(n22067), .op(n10070) );
  mux2_1 U19771 ( .ip1(\pipeline/reg_to_wr_WB [2]), .ip2(\pipeline/inst_DX [9]), .s(n22067), .op(n10068) );
  mux2_1 U19772 ( .ip1(\pipeline/reg_to_wr_WB [1]), .ip2(\pipeline/inst_DX [8]), .s(n22067), .op(n10069) );
  mux2_1 U19773 ( .ip1(\pipeline/reg_to_wr_WB [4]), .ip2(
        \pipeline/inst_DX [11]), .s(n22067), .op(n10071) );
  mux2_1 U19774 ( .ip1(\pipeline/reg_to_wr_WB [3]), .ip2(
        \pipeline/inst_DX [10]), .s(n22067), .op(n10067) );
  nand2_1 U19775 ( .ip1(\pipeline/ctrl/wr_reg_unkilled_WB ), .ip2(n22043), 
        .op(n17894) );
  nand2_1 U19776 ( .ip1(n17884), .ip2(n17883), .op(n17885) );
  nand2_1 U19777 ( .ip1(n17886), .ip2(n17885), .op(n17890) );
  nor2_1 U19778 ( .ip1(\pipeline/inst_DX [5]), .ip2(n17887), .op(n17889) );
  not_ab_or_c_or_d U19779 ( .ip1(n17891), .ip2(n17890), .ip3(n17889), .ip4(
        n17888), .op(n17892) );
  or2_1 U19780 ( .ip1(n17892), .ip2(n19505), .op(n17893) );
  nand2_1 U19781 ( .ip1(n17894), .ip2(n17893), .op(n8495) );
  nand2_1 U19782 ( .ip1(\pipeline/wb_src_sel_WB [0]), .ip2(n17895), .op(n21583) );
  nor3_1 U19783 ( .ip1(\pipeline/alu_out_WB [0]), .ip2(
        \pipeline/alu_out_WB [1]), .ip3(n21583), .op(n21238) );
  inv_1 U19784 ( .ip(\pipeline/alu_out_WB [1]), .op(n18041) );
  nor2_1 U19785 ( .ip1(n18041), .ip2(n21583), .op(n18032) );
  nand2_1 U19786 ( .ip1(\pipeline/alu_out_WB [0]), .ip2(n18032), .op(n21233)
         );
  inv_1 U19787 ( .ip(dmem_rdata[27]), .op(n17896) );
  nor2_1 U19788 ( .ip1(n21233), .ip2(n17896), .op(n17899) );
  inv_1 U19789 ( .ip(n21583), .op(n19404) );
  nand3_1 U19790 ( .ip1(\pipeline/alu_out_WB [0]), .ip2(n19404), .ip3(n18041), 
        .op(n21235) );
  inv_1 U19791 ( .ip(dmem_rdata[11]), .op(n17897) );
  nor2_1 U19792 ( .ip1(n21235), .ip2(n17897), .op(n17898) );
  not_ab_or_c_or_d U19793 ( .ip1(n21238), .ip2(dmem_rdata[3]), .ip3(n17899), 
        .ip4(n17898), .op(n17904) );
  nand2_1 U19794 ( .ip1(n17900), .ip2(n21583), .op(n17903) );
  inv_1 U19795 ( .ip(n18032), .op(n17901) );
  nor2_1 U19796 ( .ip1(\pipeline/alu_out_WB [0]), .ip2(n17901), .op(n21240) );
  nand2_1 U19797 ( .ip1(dmem_rdata[19]), .ip2(n21240), .op(n17902) );
  nand3_1 U19798 ( .ip1(n17904), .ip2(n17903), .ip3(n17902), .op(n17926) );
  nand3_1 U19799 ( .ip1(n17907), .ip2(\pipeline/reg_to_wr_WB [4]), .ip3(
        \pipeline/reg_to_wr_WB [3]), .op(n17917) );
  inv_1 U19800 ( .ip(\pipeline/reg_to_wr_WB [1]), .op(n17912) );
  nand3_1 U19801 ( .ip1(\pipeline/reg_to_wr_WB [0]), .ip2(
        \pipeline/reg_to_wr_WB [2]), .ip3(n17912), .op(n17916) );
  nor2_1 U19802 ( .ip1(n17917), .ip2(n17916), .op(n21619) );
  mux2_1 U19803 ( .ip1(\pipeline/regfile/data[29][3] ), .ip2(n17926), .s(
        n21619), .op(n8997) );
  nand3_1 U19804 ( .ip1(n17907), .ip2(\pipeline/reg_to_wr_WB [3]), .ip3(n17906), .op(n17918) );
  nand3_1 U19805 ( .ip1(\pipeline/reg_to_wr_WB [2]), .ip2(
        \pipeline/reg_to_wr_WB [1]), .ip3(n17908), .op(n17911) );
  nor2_1 U19806 ( .ip1(n17918), .ip2(n17911), .op(n21604) );
  mux2_1 U19807 ( .ip1(\pipeline/regfile/data[14][3] ), .ip2(n17926), .s(
        n21604), .op(n9477) );
  inv_1 U19808 ( .ip(\pipeline/reg_to_wr_WB [3]), .op(n17905) );
  nand3_1 U19809 ( .ip1(n17907), .ip2(\pipeline/reg_to_wr_WB [4]), .ip3(n17905), .op(n17920) );
  nor2_1 U19810 ( .ip1(n17911), .ip2(n17920), .op(n21589) );
  mux2_1 U19811 ( .ip1(\pipeline/regfile/data[22][3] ), .ip2(n17926), .s(
        n21589), .op(n9221) );
  nand3_1 U19812 ( .ip1(n17907), .ip2(n17906), .ip3(n17905), .op(n17925) );
  nor2_1 U19813 ( .ip1(n17916), .ip2(n17925), .op(n21598) );
  mux2_1 U19814 ( .ip1(\pipeline/regfile/data[5][3] ), .ip2(n17926), .s(n21598), .op(n9765) );
  nand2_1 U19815 ( .ip1(\pipeline/reg_to_wr_WB [0]), .ip2(
        \pipeline/reg_to_wr_WB [1]), .op(n17909) );
  or2_1 U19816 ( .ip1(\pipeline/reg_to_wr_WB [2]), .ip2(n17909), .op(n17921)
         );
  nor2_1 U19817 ( .ip1(n17917), .ip2(n17921), .op(n21612) );
  mux2_1 U19818 ( .ip1(\pipeline/regfile/data[27][3] ), .ip2(n17926), .s(
        n21612), .op(n9061) );
  inv_1 U19819 ( .ip(\pipeline/reg_to_wr_WB [2]), .op(n17913) );
  nand3_1 U19820 ( .ip1(\pipeline/reg_to_wr_WB [1]), .ip2(n17908), .ip3(n17913), .op(n17923) );
  nor2_1 U19821 ( .ip1(n17917), .ip2(n17923), .op(n21607) );
  mux2_1 U19822 ( .ip1(\pipeline/regfile/data[26][3] ), .ip2(n17926), .s(
        n21607), .op(n9093) );
  nor2_1 U19823 ( .ip1(\pipeline/reg_to_wr_WB [0]), .ip2(
        \pipeline/reg_to_wr_WB [1]), .op(n17914) );
  nand2_1 U19824 ( .ip1(\pipeline/reg_to_wr_WB [2]), .ip2(n17914), .op(n17924)
         );
  nor2_1 U19825 ( .ip1(n17917), .ip2(n17924), .op(n21590) );
  mux2_1 U19826 ( .ip1(\pipeline/regfile/data[28][3] ), .ip2(n17926), .s(
        n21590), .op(n9029) );
  inv_1 U19827 ( .ip(n17909), .op(n17910) );
  nand2_1 U19828 ( .ip1(\pipeline/reg_to_wr_WB [2]), .ip2(n17910), .op(n17915)
         );
  nor2_1 U19829 ( .ip1(n17917), .ip2(n17915), .op(n21606) );
  mux2_1 U19830 ( .ip1(\pipeline/regfile/data[31][3] ), .ip2(n17926), .s(
        n21606), .op(n8933) );
  nor2_1 U19831 ( .ip1(n17920), .ip2(n17921), .op(n21592) );
  mux2_1 U19832 ( .ip1(\pipeline/regfile/data[19][3] ), .ip2(n17926), .s(
        n21592), .op(n9317) );
  nor2_1 U19833 ( .ip1(n17911), .ip2(n17925), .op(n21597) );
  mux2_1 U19834 ( .ip1(\pipeline/regfile/data[6][3] ), .ip2(n17926), .s(n21597), .op(n9733) );
  nor2_1 U19835 ( .ip1(n17917), .ip2(n17911), .op(n21594) );
  mux2_1 U19836 ( .ip1(\pipeline/regfile/data[30][3] ), .ip2(n17926), .s(
        n21594), .op(n8965) );
  nor2_1 U19837 ( .ip1(n17920), .ip2(n17923), .op(n21595) );
  mux2_1 U19838 ( .ip1(\pipeline/regfile/data[18][3] ), .ip2(n17926), .s(
        n21595), .op(n9349) );
  nor2_1 U19839 ( .ip1(n17918), .ip2(n17921), .op(n21593) );
  mux2_1 U19840 ( .ip1(\pipeline/regfile/data[11][3] ), .ip2(n17926), .s(
        n21593), .op(n9573) );
  nand3_1 U19841 ( .ip1(\pipeline/reg_to_wr_WB [0]), .ip2(n17912), .ip3(n17913), .op(n17922) );
  nor2_1 U19842 ( .ip1(n17917), .ip2(n17922), .op(n21602) );
  mux2_1 U19843 ( .ip1(\pipeline/regfile/data[25][3] ), .ip2(n17926), .s(
        n21602), .op(n9125) );
  nor2_1 U19844 ( .ip1(n17916), .ip2(n17918), .op(n21600) );
  mux2_1 U19845 ( .ip1(\pipeline/regfile/data[13][3] ), .ip2(n17926), .s(
        n21600), .op(n9509) );
  nor2_1 U19846 ( .ip1(n17920), .ip2(n17922), .op(n21616) );
  mux2_1 U19847 ( .ip1(\pipeline/regfile/data[17][3] ), .ip2(n17926), .s(
        n21616), .op(n9381) );
  nor2_1 U19848 ( .ip1(n17920), .ip2(n17915), .op(n21596) );
  mux2_1 U19849 ( .ip1(\pipeline/regfile/data[23][3] ), .ip2(n17926), .s(
        n21596), .op(n9189) );
  nor2_1 U19850 ( .ip1(n17918), .ip2(n17924), .op(n21591) );
  mux2_1 U19851 ( .ip1(\pipeline/regfile/data[12][3] ), .ip2(n17926), .s(
        n21591), .op(n9541) );
  nor2_1 U19852 ( .ip1(n17925), .ip2(n17915), .op(n21614) );
  mux2_1 U19853 ( .ip1(\pipeline/regfile/data[7][3] ), .ip2(n17926), .s(n21614), .op(n9701) );
  nand2_1 U19854 ( .ip1(n17914), .ip2(n17913), .op(n17919) );
  nor2_1 U19855 ( .ip1(n17918), .ip2(n17919), .op(n21617) );
  mux2_1 U19856 ( .ip1(\pipeline/regfile/data[8][3] ), .ip2(n17926), .s(n21617), .op(n9669) );
  nor2_1 U19857 ( .ip1(n17918), .ip2(n17915), .op(n21613) );
  mux2_1 U19858 ( .ip1(\pipeline/regfile/data[15][3] ), .ip2(n17926), .s(
        n21613), .op(n9445) );
  nor2_1 U19859 ( .ip1(n17918), .ip2(n17923), .op(n21618) );
  mux2_1 U19860 ( .ip1(\pipeline/regfile/data[10][3] ), .ip2(n17926), .s(
        n21618), .op(n9605) );
  nor2_1 U19861 ( .ip1(n17916), .ip2(n17920), .op(n21615) );
  mux2_1 U19862 ( .ip1(\pipeline/regfile/data[21][3] ), .ip2(n17926), .s(
        n21615), .op(n9253) );
  nor2_1 U19863 ( .ip1(n17917), .ip2(n17919), .op(n21603) );
  mux2_1 U19864 ( .ip1(\pipeline/regfile/data[24][3] ), .ip2(n17926), .s(
        n21603), .op(n9157) );
  nor2_1 U19865 ( .ip1(n17920), .ip2(n17924), .op(n21601) );
  mux2_1 U19866 ( .ip1(\pipeline/regfile/data[20][3] ), .ip2(n17926), .s(
        n21601), .op(n9285) );
  nor2_1 U19867 ( .ip1(n17918), .ip2(n17922), .op(n21609) );
  mux2_1 U19868 ( .ip1(\pipeline/regfile/data[9][3] ), .ip2(n17926), .s(n21609), .op(n9637) );
  nor2_1 U19869 ( .ip1(n17920), .ip2(n17919), .op(n21608) );
  mux2_1 U19870 ( .ip1(\pipeline/regfile/data[16][3] ), .ip2(n17926), .s(
        n21608), .op(n9413) );
  nor2_1 U19871 ( .ip1(n17925), .ip2(n17921), .op(n21599) );
  mux2_1 U19872 ( .ip1(\pipeline/regfile/data[3][3] ), .ip2(n17926), .s(n21599), .op(n9829) );
  nor2_1 U19873 ( .ip1(n17925), .ip2(n17922), .op(n21611) );
  mux2_1 U19874 ( .ip1(\pipeline/regfile/data[1][3] ), .ip2(n17926), .s(n21611), .op(n9893) );
  nor2_1 U19875 ( .ip1(n17925), .ip2(n17923), .op(n21610) );
  mux2_1 U19876 ( .ip1(\pipeline/regfile/data[2][3] ), .ip2(n17926), .s(n21610), .op(n9861) );
  nor2_1 U19877 ( .ip1(n17925), .ip2(n17924), .op(n21605) );
  mux2_1 U19878 ( .ip1(\pipeline/regfile/data[4][3] ), .ip2(n17926), .s(n21605), .op(n9797) );
  inv_1 U19879 ( .ip(dmem_rdata[28]), .op(n17927) );
  nor2_1 U19880 ( .ip1(n21233), .ip2(n17927), .op(n17930) );
  inv_1 U19881 ( .ip(dmem_rdata[12]), .op(n17928) );
  nor2_1 U19882 ( .ip1(n21235), .ip2(n17928), .op(n17929) );
  not_ab_or_c_or_d U19883 ( .ip1(n21238), .ip2(dmem_rdata[4]), .ip3(n17930), 
        .ip4(n17929), .op(n17934) );
  nand2_1 U19884 ( .ip1(n17931), .ip2(n21583), .op(n17933) );
  nand2_1 U19885 ( .ip1(n21240), .ip2(dmem_rdata[20]), .op(n17932) );
  nand3_1 U19886 ( .ip1(n17934), .ip2(n17933), .ip3(n17932), .op(n17935) );
  mux2_1 U19887 ( .ip1(\pipeline/regfile/data[22][4] ), .ip2(n17935), .s(
        n21589), .op(n9220) );
  mux2_1 U19888 ( .ip1(\pipeline/regfile/data[28][4] ), .ip2(n17935), .s(
        n21590), .op(n9028) );
  mux2_1 U19889 ( .ip1(\pipeline/regfile/data[12][4] ), .ip2(n17935), .s(
        n21591), .op(n9540) );
  mux2_1 U19890 ( .ip1(\pipeline/regfile/data[19][4] ), .ip2(n17935), .s(
        n21592), .op(n9316) );
  mux2_1 U19891 ( .ip1(\pipeline/regfile/data[11][4] ), .ip2(n17935), .s(
        n21593), .op(n9572) );
  mux2_1 U19892 ( .ip1(\pipeline/regfile/data[30][4] ), .ip2(n17935), .s(
        n21594), .op(n8964) );
  mux2_1 U19893 ( .ip1(\pipeline/regfile/data[18][4] ), .ip2(n17935), .s(
        n21595), .op(n9348) );
  mux2_1 U19894 ( .ip1(\pipeline/regfile/data[23][4] ), .ip2(n17935), .s(
        n21596), .op(n9188) );
  mux2_1 U19895 ( .ip1(\pipeline/regfile/data[6][4] ), .ip2(n17935), .s(n21597), .op(n9732) );
  mux2_1 U19896 ( .ip1(\pipeline/regfile/data[5][4] ), .ip2(n17935), .s(n21598), .op(n9764) );
  mux2_1 U19897 ( .ip1(\pipeline/regfile/data[3][4] ), .ip2(n17935), .s(n21599), .op(n9828) );
  mux2_1 U19898 ( .ip1(\pipeline/regfile/data[13][4] ), .ip2(n17935), .s(
        n21600), .op(n9508) );
  mux2_1 U19899 ( .ip1(\pipeline/regfile/data[20][4] ), .ip2(n17935), .s(
        n21601), .op(n9284) );
  mux2_1 U19900 ( .ip1(\pipeline/regfile/data[25][4] ), .ip2(n17935), .s(
        n21602), .op(n9124) );
  mux2_1 U19901 ( .ip1(\pipeline/regfile/data[24][4] ), .ip2(n17935), .s(
        n21603), .op(n9156) );
  mux2_1 U19902 ( .ip1(\pipeline/regfile/data[14][4] ), .ip2(n17935), .s(
        n21604), .op(n9476) );
  mux2_1 U19903 ( .ip1(\pipeline/regfile/data[4][4] ), .ip2(n17935), .s(n21605), .op(n9796) );
  mux2_1 U19904 ( .ip1(\pipeline/regfile/data[31][4] ), .ip2(n17935), .s(
        n21606), .op(n8932) );
  mux2_1 U19905 ( .ip1(\pipeline/regfile/data[26][4] ), .ip2(n17935), .s(
        n21607), .op(n9092) );
  mux2_1 U19906 ( .ip1(\pipeline/regfile/data[16][4] ), .ip2(n17935), .s(
        n21608), .op(n9412) );
  mux2_1 U19907 ( .ip1(\pipeline/regfile/data[9][4] ), .ip2(n17935), .s(n21609), .op(n9636) );
  mux2_1 U19908 ( .ip1(\pipeline/regfile/data[2][4] ), .ip2(n17935), .s(n21610), .op(n9860) );
  mux2_1 U19909 ( .ip1(\pipeline/regfile/data[1][4] ), .ip2(n17935), .s(n21611), .op(n9892) );
  mux2_1 U19910 ( .ip1(\pipeline/regfile/data[27][4] ), .ip2(n17935), .s(
        n21612), .op(n9060) );
  mux2_1 U19911 ( .ip1(\pipeline/regfile/data[15][4] ), .ip2(n17935), .s(
        n21613), .op(n9444) );
  mux2_1 U19912 ( .ip1(\pipeline/regfile/data[7][4] ), .ip2(n17935), .s(n21614), .op(n9700) );
  mux2_1 U19913 ( .ip1(\pipeline/regfile/data[21][4] ), .ip2(n17935), .s(
        n21615), .op(n9252) );
  mux2_1 U19914 ( .ip1(\pipeline/regfile/data[17][4] ), .ip2(n17935), .s(
        n21616), .op(n9380) );
  mux2_1 U19915 ( .ip1(\pipeline/regfile/data[8][4] ), .ip2(n17935), .s(n21617), .op(n9668) );
  mux2_1 U19916 ( .ip1(\pipeline/regfile/data[10][4] ), .ip2(n17935), .s(
        n21618), .op(n9604) );
  mux2_1 U19917 ( .ip1(\pipeline/regfile/data[29][4] ), .ip2(n17935), .s(
        n21619), .op(n8996) );
  nand2_1 U19918 ( .ip1(n19498), .ip2(dmem_htrans[1]), .op(n17937) );
  nand2_1 U19919 ( .ip1(\pipeline/ctrl/dmem_en_WB ), .ip2(n22043), .op(n17936)
         );
  nand2_1 U19920 ( .ip1(n17937), .ip2(n17936), .op(n8497) );
  nor2_1 U19921 ( .ip1(n17938), .ip2(n20483), .op(n17940) );
  xor2_1 U19922 ( .ip1(n17940), .ip2(n17939), .op(n17941) );
  nand2_1 U19923 ( .ip1(n21649), .ip2(n17941), .op(n17947) );
  nor3_1 U19924 ( .ip1(n21884), .ip2(n17943), .ip3(n17942), .op(n17944) );
  xor2_1 U19925 ( .ip1(\pipeline/md/a [4]), .ip2(n17944), .op(n17945) );
  nand2_1 U19926 ( .ip1(n14770), .ip2(n22665), .op(n21643) );
  nand2_1 U19927 ( .ip1(n17945), .ip2(n21643), .op(n17946) );
  nand2_1 U19928 ( .ip1(n17947), .ip2(n17946), .op(n8390) );
  nand2_1 U19929 ( .ip1(n17949), .ip2(n17948), .op(n17950) );
  nand2_1 U19930 ( .ip1(n17951), .ip2(n17950), .op(n22360) );
  nor2_1 U19931 ( .ip1(n21029), .ip2(n22360), .op(n17955) );
  inv_1 U19932 ( .ip(\pipeline/csr/mtvec [4]), .op(n17952) );
  nor2_1 U19933 ( .ip1(htif_reset), .ip2(n17952), .op(n17953) );
  nor2_1 U19934 ( .ip1(n21032), .ip2(n17953), .op(n17954) );
  nor2_1 U19935 ( .ip1(n17955), .ip2(n17954), .op(n9988) );
  xor2_1 U19936 ( .ip1(n17957), .ip2(n17956), .op(n17961) );
  inv_1 U19937 ( .ip(n21161), .op(n17958) );
  nand2_1 U19938 ( .ip1(n21162), .ip2(n17958), .op(n17959) );
  nand2_1 U19939 ( .ip1(n17959), .ip2(n14208), .op(n17960) );
  xor2_1 U19940 ( .ip1(n17961), .ip2(n17960), .op(imem_haddr[4]) );
  nand2_1 U19941 ( .ip1(n21995), .ip2(imem_haddr[4]), .op(n17963) );
  nand2_1 U19942 ( .ip1(\pipeline/PC_IF [4]), .ip2(n21996), .op(n17962) );
  nand2_1 U19943 ( .ip1(n17963), .ip2(n17962), .op(n8482) );
  nand2_1 U19944 ( .ip1(\pipeline/PC_IF [4]), .ip2(n21988), .op(n17965) );
  nand2_1 U19945 ( .ip1(\pipeline/PC_DX [4]), .ip2(n21999), .op(n17964) );
  nand2_1 U19946 ( .ip1(n17965), .ip2(n17964), .op(n8481) );
  mux2_1 U19947 ( .ip1(\pipeline/PC_WB [4]), .ip2(\pipeline/PC_DX [4]), .s(
        n22067), .op(n8899) );
  inv_1 U19948 ( .ip(n21174), .op(n18637) );
  nor2_1 U19949 ( .ip1(n17966), .ip2(n18637), .op(n17971) );
  inv_1 U19950 ( .ip(\pipeline/PC_WB [4]), .op(n17969) );
  inv_1 U19951 ( .ip(n21169), .op(n17967) );
  nand2_1 U19952 ( .ip1(n17967), .ip2(\pipeline/PC_WB [3]), .op(n17968) );
  not_ab_or_c_or_d U19953 ( .ip1(n17969), .ip2(n17968), .ip3(n21044), .ip4(
        n21171), .op(n17970) );
  ab_or_c_or_d U19954 ( .ip1(n21043), .ip2(n17972), .ip3(n17971), .ip4(n17970), 
        .op(n8867) );
  mux2_1 U19955 ( .ip1(\pipeline/PC_WB [12]), .ip2(\pipeline/PC_DX [12]), .s(
        n20389), .op(n8891) );
  mux2_1 U19956 ( .ip1(\pipeline/csr_rdata_WB [5]), .ip2(n17973), .s(n19498), 
        .op(n8801) );
  inv_1 U19957 ( .ip(dmem_rdata[29]), .op(n17974) );
  nor2_1 U19958 ( .ip1(n21233), .ip2(n17974), .op(n17977) );
  inv_1 U19959 ( .ip(dmem_rdata[13]), .op(n17975) );
  nor2_1 U19960 ( .ip1(n21235), .ip2(n17975), .op(n17976) );
  not_ab_or_c_or_d U19961 ( .ip1(n21238), .ip2(dmem_rdata[5]), .ip3(n17977), 
        .ip4(n17976), .op(n17981) );
  nand2_1 U19962 ( .ip1(n17978), .ip2(n21583), .op(n17980) );
  nand2_1 U19963 ( .ip1(n21240), .ip2(dmem_rdata[21]), .op(n17979) );
  nand3_1 U19964 ( .ip1(n17981), .ip2(n17980), .ip3(n17979), .op(n17982) );
  mux2_1 U19965 ( .ip1(\pipeline/regfile/data[29][5] ), .ip2(n17982), .s(
        n21619), .op(n8995) );
  mux2_1 U19966 ( .ip1(\pipeline/regfile/data[14][5] ), .ip2(n17982), .s(
        n21604), .op(n9475) );
  mux2_1 U19967 ( .ip1(\pipeline/regfile/data[22][5] ), .ip2(n17982), .s(
        n21589), .op(n9219) );
  mux2_1 U19968 ( .ip1(\pipeline/regfile/data[5][5] ), .ip2(n17982), .s(n21598), .op(n9763) );
  mux2_1 U19969 ( .ip1(\pipeline/regfile/data[27][5] ), .ip2(n17982), .s(
        n21612), .op(n9059) );
  mux2_1 U19970 ( .ip1(\pipeline/regfile/data[26][5] ), .ip2(n17982), .s(
        n21607), .op(n9091) );
  mux2_1 U19971 ( .ip1(\pipeline/regfile/data[28][5] ), .ip2(n17982), .s(
        n21590), .op(n9027) );
  mux2_1 U19972 ( .ip1(\pipeline/regfile/data[31][5] ), .ip2(n17982), .s(
        n21606), .op(n8931) );
  mux2_1 U19973 ( .ip1(\pipeline/regfile/data[19][5] ), .ip2(n17982), .s(
        n21592), .op(n9315) );
  mux2_1 U19974 ( .ip1(\pipeline/regfile/data[6][5] ), .ip2(n17982), .s(n21597), .op(n9731) );
  mux2_1 U19975 ( .ip1(\pipeline/regfile/data[30][5] ), .ip2(n17982), .s(
        n21594), .op(n8963) );
  mux2_1 U19976 ( .ip1(\pipeline/regfile/data[18][5] ), .ip2(n17982), .s(
        n21595), .op(n9347) );
  mux2_1 U19977 ( .ip1(\pipeline/regfile/data[11][5] ), .ip2(n17982), .s(
        n21593), .op(n9571) );
  mux2_1 U19978 ( .ip1(\pipeline/regfile/data[25][5] ), .ip2(n17982), .s(
        n21602), .op(n9123) );
  mux2_1 U19979 ( .ip1(\pipeline/regfile/data[13][5] ), .ip2(n17982), .s(
        n21600), .op(n9507) );
  mux2_1 U19980 ( .ip1(\pipeline/regfile/data[17][5] ), .ip2(n17982), .s(
        n21616), .op(n9379) );
  mux2_1 U19981 ( .ip1(\pipeline/regfile/data[23][5] ), .ip2(n17982), .s(
        n21596), .op(n9187) );
  mux2_1 U19982 ( .ip1(\pipeline/regfile/data[12][5] ), .ip2(n17982), .s(
        n21591), .op(n9539) );
  mux2_1 U19983 ( .ip1(\pipeline/regfile/data[7][5] ), .ip2(n17982), .s(n21614), .op(n9699) );
  mux2_1 U19984 ( .ip1(\pipeline/regfile/data[8][5] ), .ip2(n17982), .s(n21617), .op(n9667) );
  mux2_1 U19985 ( .ip1(\pipeline/regfile/data[15][5] ), .ip2(n17982), .s(
        n21613), .op(n9443) );
  mux2_1 U19986 ( .ip1(\pipeline/regfile/data[10][5] ), .ip2(n17982), .s(
        n21618), .op(n9603) );
  mux2_1 U19987 ( .ip1(\pipeline/regfile/data[21][5] ), .ip2(n17982), .s(
        n21615), .op(n9251) );
  mux2_1 U19988 ( .ip1(\pipeline/regfile/data[24][5] ), .ip2(n17982), .s(
        n21603), .op(n9155) );
  mux2_1 U19989 ( .ip1(\pipeline/regfile/data[20][5] ), .ip2(n17982), .s(
        n21601), .op(n9283) );
  mux2_1 U19990 ( .ip1(\pipeline/regfile/data[9][5] ), .ip2(n17982), .s(n21609), .op(n9635) );
  mux2_1 U19991 ( .ip1(\pipeline/regfile/data[16][5] ), .ip2(n17982), .s(
        n21608), .op(n9411) );
  mux2_1 U19992 ( .ip1(\pipeline/regfile/data[3][5] ), .ip2(n17982), .s(n21599), .op(n9827) );
  mux2_1 U19993 ( .ip1(\pipeline/regfile/data[1][5] ), .ip2(n17982), .s(n21611), .op(n9891) );
  mux2_1 U19994 ( .ip1(\pipeline/regfile/data[2][5] ), .ip2(n17982), .s(n21610), .op(n9859) );
  mux2_1 U19995 ( .ip1(\pipeline/regfile/data[4][5] ), .ip2(n17982), .s(n21605), .op(n9795) );
  nor2_1 U19996 ( .ip1(n21029), .ip2(n22364), .op(n17986) );
  inv_1 U19997 ( .ip(\pipeline/csr/mtvec [6]), .op(n17983) );
  nor2_1 U19998 ( .ip1(htif_reset), .ip2(n17983), .op(n17984) );
  nor2_1 U19999 ( .ip1(n21032), .ip2(n17984), .op(n17985) );
  nor2_1 U20000 ( .ip1(n17986), .ip2(n17985), .op(n9986) );
  nor2_1 U20001 ( .ip1(n18229), .ip2(n18232), .op(n17993) );
  inv_1 U20002 ( .ip(n17987), .op(n17988) );
  nand2_1 U20003 ( .ip1(n17989), .ip2(n17988), .op(n21037) );
  inv_1 U20004 ( .ip(n21036), .op(n17990) );
  nand2_1 U20005 ( .ip1(n21037), .ip2(n17990), .op(n17992) );
  inv_1 U20006 ( .ip(n21035), .op(n17991) );
  nand2_1 U20007 ( .ip1(n17992), .ip2(n17991), .op(n18231) );
  xor2_1 U20008 ( .ip1(n17993), .ip2(n18231), .op(imem_haddr[6]) );
  nand2_1 U20009 ( .ip1(n21995), .ip2(imem_haddr[6]), .op(n17995) );
  nand2_1 U20010 ( .ip1(\pipeline/PC_IF [6]), .ip2(n21996), .op(n17994) );
  nand2_1 U20011 ( .ip1(n17995), .ip2(n17994), .op(n8478) );
  nand2_1 U20012 ( .ip1(\pipeline/PC_IF [6]), .ip2(n21988), .op(n17997) );
  nand2_1 U20013 ( .ip1(\pipeline/PC_DX [6]), .ip2(n21999), .op(n17996) );
  nand2_1 U20014 ( .ip1(n17997), .ip2(n17996), .op(n8477) );
  mux2_1 U20015 ( .ip1(\pipeline/PC_WB [6]), .ip2(\pipeline/PC_DX [6]), .s(
        n22067), .op(n8897) );
  nand2_1 U20016 ( .ip1(n21043), .ip2(n22364), .op(n18002) );
  inv_1 U20017 ( .ip(n17998), .op(n19681) );
  xor2_1 U20018 ( .ip1(n19681), .ip2(\pipeline/PC_WB [6]), .op(n17999) );
  nand2_1 U20019 ( .ip1(n21046), .ip2(n17999), .op(n18001) );
  nand2_1 U20020 ( .ip1(\pipeline/epc [6]), .ip2(n21174), .op(n18000) );
  nand3_1 U20021 ( .ip1(n18002), .ip2(n18001), .ip3(n18000), .op(n8865) );
  inv_1 U20022 ( .ip(dmem_rdata[30]), .op(n18003) );
  nor2_1 U20023 ( .ip1(n21233), .ip2(n18003), .op(n18006) );
  inv_1 U20024 ( .ip(dmem_rdata[14]), .op(n18004) );
  nor2_1 U20025 ( .ip1(n21235), .ip2(n18004), .op(n18005) );
  not_ab_or_c_or_d U20026 ( .ip1(n21238), .ip2(dmem_rdata[6]), .ip3(n18006), 
        .ip4(n18005), .op(n18010) );
  nand2_1 U20027 ( .ip1(n18007), .ip2(n21583), .op(n18009) );
  nand2_1 U20028 ( .ip1(n21240), .ip2(dmem_rdata[22]), .op(n18008) );
  nand3_1 U20029 ( .ip1(n18010), .ip2(n18009), .ip3(n18008), .op(n18011) );
  mux2_1 U20030 ( .ip1(\pipeline/regfile/data[29][6] ), .ip2(n18011), .s(
        n21619), .op(n8994) );
  mux2_1 U20031 ( .ip1(\pipeline/regfile/data[14][6] ), .ip2(n18011), .s(
        n21604), .op(n9474) );
  mux2_1 U20032 ( .ip1(\pipeline/regfile/data[22][6] ), .ip2(n18011), .s(
        n21589), .op(n9218) );
  mux2_1 U20033 ( .ip1(\pipeline/regfile/data[5][6] ), .ip2(n18011), .s(n21598), .op(n9762) );
  mux2_1 U20034 ( .ip1(\pipeline/regfile/data[27][6] ), .ip2(n18011), .s(
        n21612), .op(n9058) );
  mux2_1 U20035 ( .ip1(\pipeline/regfile/data[26][6] ), .ip2(n18011), .s(
        n21607), .op(n9090) );
  mux2_1 U20036 ( .ip1(\pipeline/regfile/data[28][6] ), .ip2(n18011), .s(
        n21590), .op(n9026) );
  mux2_1 U20037 ( .ip1(\pipeline/regfile/data[31][6] ), .ip2(n18011), .s(
        n21606), .op(n8930) );
  mux2_1 U20038 ( .ip1(\pipeline/regfile/data[19][6] ), .ip2(n18011), .s(
        n21592), .op(n9314) );
  mux2_1 U20039 ( .ip1(\pipeline/regfile/data[6][6] ), .ip2(n18011), .s(n21597), .op(n9730) );
  mux2_1 U20040 ( .ip1(\pipeline/regfile/data[30][6] ), .ip2(n18011), .s(
        n21594), .op(n8962) );
  mux2_1 U20041 ( .ip1(\pipeline/regfile/data[18][6] ), .ip2(n18011), .s(
        n21595), .op(n9346) );
  mux2_1 U20042 ( .ip1(\pipeline/regfile/data[11][6] ), .ip2(n18011), .s(
        n21593), .op(n9570) );
  mux2_1 U20043 ( .ip1(\pipeline/regfile/data[25][6] ), .ip2(n18011), .s(
        n21602), .op(n9122) );
  mux2_1 U20044 ( .ip1(\pipeline/regfile/data[13][6] ), .ip2(n18011), .s(
        n21600), .op(n9506) );
  mux2_1 U20045 ( .ip1(\pipeline/regfile/data[17][6] ), .ip2(n18011), .s(
        n21616), .op(n9378) );
  mux2_1 U20046 ( .ip1(\pipeline/regfile/data[23][6] ), .ip2(n18011), .s(
        n21596), .op(n9186) );
  mux2_1 U20047 ( .ip1(\pipeline/regfile/data[12][6] ), .ip2(n18011), .s(
        n21591), .op(n9538) );
  mux2_1 U20048 ( .ip1(\pipeline/regfile/data[7][6] ), .ip2(n18011), .s(n21614), .op(n9698) );
  mux2_1 U20049 ( .ip1(\pipeline/regfile/data[8][6] ), .ip2(n18011), .s(n21617), .op(n9666) );
  mux2_1 U20050 ( .ip1(\pipeline/regfile/data[15][6] ), .ip2(n18011), .s(
        n21613), .op(n9442) );
  mux2_1 U20051 ( .ip1(\pipeline/regfile/data[10][6] ), .ip2(n18011), .s(
        n21618), .op(n9602) );
  mux2_1 U20052 ( .ip1(\pipeline/regfile/data[21][6] ), .ip2(n18011), .s(
        n21615), .op(n9250) );
  mux2_1 U20053 ( .ip1(\pipeline/regfile/data[24][6] ), .ip2(n18011), .s(
        n21603), .op(n9154) );
  mux2_1 U20054 ( .ip1(\pipeline/regfile/data[20][6] ), .ip2(n18011), .s(
        n21601), .op(n9282) );
  mux2_1 U20055 ( .ip1(\pipeline/regfile/data[9][6] ), .ip2(n18011), .s(n21609), .op(n9634) );
  mux2_1 U20056 ( .ip1(\pipeline/regfile/data[16][6] ), .ip2(n18011), .s(
        n21608), .op(n9410) );
  mux2_1 U20057 ( .ip1(\pipeline/regfile/data[3][6] ), .ip2(n18011), .s(n21599), .op(n9826) );
  mux2_1 U20058 ( .ip1(\pipeline/regfile/data[1][6] ), .ip2(n18011), .s(n21611), .op(n9890) );
  mux2_1 U20059 ( .ip1(\pipeline/regfile/data[2][6] ), .ip2(n18011), .s(n21610), .op(n9858) );
  mux2_1 U20060 ( .ip1(\pipeline/regfile/data[4][6] ), .ip2(n18011), .s(n21605), .op(n9794) );
  inv_1 U20061 ( .ip(dmem_rdata[25]), .op(n18012) );
  nor2_1 U20062 ( .ip1(n21233), .ip2(n18012), .op(n18015) );
  inv_1 U20063 ( .ip(dmem_rdata[9]), .op(n18013) );
  nor2_1 U20064 ( .ip1(n21235), .ip2(n18013), .op(n18014) );
  not_ab_or_c_or_d U20065 ( .ip1(n21238), .ip2(dmem_rdata[1]), .ip3(n18015), 
        .ip4(n18014), .op(n18019) );
  nand2_1 U20066 ( .ip1(n18016), .ip2(n21583), .op(n18018) );
  nand2_1 U20067 ( .ip1(n21240), .ip2(dmem_rdata[17]), .op(n18017) );
  nand3_1 U20068 ( .ip1(n18019), .ip2(n18018), .ip3(n18017), .op(n18020) );
  mux2_1 U20069 ( .ip1(\pipeline/regfile/data[22][1] ), .ip2(n18020), .s(
        n21589), .op(n9223) );
  mux2_1 U20070 ( .ip1(\pipeline/regfile/data[28][1] ), .ip2(n18020), .s(
        n21590), .op(n9031) );
  mux2_1 U20071 ( .ip1(\pipeline/regfile/data[12][1] ), .ip2(n18020), .s(
        n21591), .op(n9543) );
  mux2_1 U20072 ( .ip1(\pipeline/regfile/data[19][1] ), .ip2(n18020), .s(
        n21592), .op(n9319) );
  mux2_1 U20073 ( .ip1(\pipeline/regfile/data[11][1] ), .ip2(n18020), .s(
        n21593), .op(n9575) );
  mux2_1 U20074 ( .ip1(\pipeline/regfile/data[30][1] ), .ip2(n18020), .s(
        n21594), .op(n8967) );
  mux2_1 U20075 ( .ip1(\pipeline/regfile/data[18][1] ), .ip2(n18020), .s(
        n21595), .op(n9351) );
  mux2_1 U20076 ( .ip1(\pipeline/regfile/data[23][1] ), .ip2(n18020), .s(
        n21596), .op(n9191) );
  mux2_1 U20077 ( .ip1(\pipeline/regfile/data[6][1] ), .ip2(n18020), .s(n21597), .op(n9735) );
  mux2_1 U20078 ( .ip1(\pipeline/regfile/data[5][1] ), .ip2(n18020), .s(n21598), .op(n9767) );
  mux2_1 U20079 ( .ip1(\pipeline/regfile/data[3][1] ), .ip2(n18020), .s(n21599), .op(n9831) );
  mux2_1 U20080 ( .ip1(\pipeline/regfile/data[13][1] ), .ip2(n18020), .s(
        n21600), .op(n9511) );
  mux2_1 U20081 ( .ip1(\pipeline/regfile/data[20][1] ), .ip2(n18020), .s(
        n21601), .op(n9287) );
  mux2_1 U20082 ( .ip1(\pipeline/regfile/data[25][1] ), .ip2(n18020), .s(
        n21602), .op(n9127) );
  mux2_1 U20083 ( .ip1(\pipeline/regfile/data[24][1] ), .ip2(n18020), .s(
        n21603), .op(n9159) );
  mux2_1 U20084 ( .ip1(\pipeline/regfile/data[14][1] ), .ip2(n18020), .s(
        n21604), .op(n9479) );
  mux2_1 U20085 ( .ip1(\pipeline/regfile/data[4][1] ), .ip2(n18020), .s(n21605), .op(n9799) );
  mux2_1 U20086 ( .ip1(\pipeline/regfile/data[31][1] ), .ip2(n18020), .s(
        n21606), .op(n8935) );
  mux2_1 U20087 ( .ip1(\pipeline/regfile/data[26][1] ), .ip2(n18020), .s(
        n21607), .op(n9095) );
  mux2_1 U20088 ( .ip1(\pipeline/regfile/data[16][1] ), .ip2(n18020), .s(
        n21608), .op(n9415) );
  mux2_1 U20089 ( .ip1(\pipeline/regfile/data[9][1] ), .ip2(n18020), .s(n21609), .op(n9639) );
  mux2_1 U20090 ( .ip1(\pipeline/regfile/data[2][1] ), .ip2(n18020), .s(n21610), .op(n9863) );
  mux2_1 U20091 ( .ip1(\pipeline/regfile/data[1][1] ), .ip2(n18020), .s(n21611), .op(n9895) );
  mux2_1 U20092 ( .ip1(\pipeline/regfile/data[27][1] ), .ip2(n18020), .s(
        n21612), .op(n9063) );
  mux2_1 U20093 ( .ip1(\pipeline/regfile/data[15][1] ), .ip2(n18020), .s(
        n21613), .op(n9447) );
  mux2_1 U20094 ( .ip1(\pipeline/regfile/data[7][1] ), .ip2(n18020), .s(n21614), .op(n9703) );
  mux2_1 U20095 ( .ip1(\pipeline/regfile/data[21][1] ), .ip2(n18020), .s(
        n21615), .op(n9255) );
  mux2_1 U20096 ( .ip1(\pipeline/regfile/data[17][1] ), .ip2(n18020), .s(
        n21616), .op(n9383) );
  mux2_1 U20097 ( .ip1(\pipeline/regfile/data[8][1] ), .ip2(n18020), .s(n21617), .op(n9671) );
  mux2_1 U20098 ( .ip1(\pipeline/regfile/data[10][1] ), .ip2(n18020), .s(
        n21618), .op(n9607) );
  mux2_1 U20099 ( .ip1(\pipeline/regfile/data[29][1] ), .ip2(n18020), .s(
        n21619), .op(n8999) );
  nand2_1 U20100 ( .ip1(\pipeline/PC_DX [0]), .ip2(n18021), .op(n18027) );
  nand2_1 U20101 ( .ip1(n18023), .ip2(n18022), .op(n18026) );
  nand2_1 U20102 ( .ip1(n18024), .ip2(\pipeline/PC_IF [0]), .op(n18025) );
  nand3_1 U20103 ( .ip1(n18027), .ip2(n18026), .ip3(n18025), .op(imem_haddr[0]) );
  nand2_1 U20104 ( .ip1(n21995), .ip2(imem_haddr[0]), .op(n18029) );
  nand2_1 U20105 ( .ip1(n21996), .ip2(\pipeline/PC_IF [0]), .op(n18028) );
  nand2_1 U20106 ( .ip1(n18029), .ip2(n18028), .op(n8490) );
  nand2_1 U20107 ( .ip1(n21988), .ip2(\pipeline/PC_IF [0]), .op(n18031) );
  nand2_1 U20108 ( .ip1(\pipeline/PC_DX [0]), .ip2(n21999), .op(n18030) );
  nand2_1 U20109 ( .ip1(n18031), .ip2(n18030), .op(n8489) );
  or2_1 U20110 ( .ip1(\pipeline/dmem_type_WB [1]), .ip2(
        \pipeline/dmem_type_WB [2]), .op(n22344) );
  mux2_1 U20111 ( .ip1(dmem_rdata[23]), .ip2(dmem_rdata[31]), .s(
        \pipeline/alu_out_WB [0]), .op(n19303) );
  nand2_1 U20112 ( .ip1(n18032), .ip2(n19303), .op(n18035) );
  nand2_1 U20113 ( .ip1(n21238), .ip2(dmem_rdata[7]), .op(n18034) );
  inv_1 U20114 ( .ip(n21235), .op(n19386) );
  nand2_1 U20115 ( .ip1(n19386), .ip2(dmem_rdata[15]), .op(n18033) );
  and3_1 U20116 ( .ip1(n18035), .ip2(n18034), .ip3(n18033), .op(n18245) );
  nor3_1 U20117 ( .ip1(n22344), .ip2(\pipeline/dmem_type_WB [0]), .ip3(n18245), 
        .op(n19390) );
  mux2_1 U20118 ( .ip1(dmem_rdata[15]), .ip2(dmem_rdata[23]), .s(
        \pipeline/alu_out_WB [0]), .op(n18036) );
  inv_1 U20119 ( .ip(n18036), .op(n18038) );
  inv_1 U20120 ( .ip(\pipeline/alu_out_WB [0]), .op(n18516) );
  nand2_1 U20121 ( .ip1(dmem_rdata[31]), .ip2(n18516), .op(n18037) );
  mux2_1 U20122 ( .ip1(n18038), .ip2(n18037), .s(\pipeline/alu_out_WB [1]), 
        .op(n18281) );
  inv_1 U20123 ( .ip(n22344), .op(n22087) );
  nand2_1 U20124 ( .ip1(n22087), .ip2(\pipeline/dmem_type_WB [0]), .op(n22321)
         );
  nor3_1 U20125 ( .ip1(n21583), .ip2(n18281), .ip3(n22321), .op(n18039) );
  nor2_1 U20126 ( .ip1(n19390), .ip2(n18039), .op(n21588) );
  nand2_1 U20127 ( .ip1(n18040), .ip2(n21583), .op(n18043) );
  nand3_1 U20128 ( .ip1(\pipeline/dmem_type_WB [1]), .ip2(n19404), .ip3(n18041), .op(n19302) );
  nor2_1 U20129 ( .ip1(\pipeline/alu_out_WB [0]), .ip2(n19302), .op(n21585) );
  nand2_1 U20130 ( .ip1(dmem_rdata[29]), .ip2(n21585), .op(n18042) );
  nand3_1 U20131 ( .ip1(n21588), .ip2(n18043), .ip3(n18042), .op(n18044) );
  mux2_1 U20132 ( .ip1(\pipeline/regfile/data[22][29] ), .ip2(n18044), .s(
        n21589), .op(n9195) );
  mux2_1 U20133 ( .ip1(\pipeline/regfile/data[28][29] ), .ip2(n18044), .s(
        n21590), .op(n9003) );
  mux2_1 U20134 ( .ip1(\pipeline/regfile/data[12][29] ), .ip2(n18044), .s(
        n21591), .op(n9515) );
  mux2_1 U20135 ( .ip1(\pipeline/regfile/data[19][29] ), .ip2(n18044), .s(
        n21592), .op(n9291) );
  mux2_1 U20136 ( .ip1(\pipeline/regfile/data[11][29] ), .ip2(n18044), .s(
        n21593), .op(n9547) );
  mux2_1 U20137 ( .ip1(\pipeline/regfile/data[30][29] ), .ip2(n18044), .s(
        n21594), .op(n8939) );
  mux2_1 U20138 ( .ip1(\pipeline/regfile/data[18][29] ), .ip2(n18044), .s(
        n21595), .op(n9323) );
  mux2_1 U20139 ( .ip1(\pipeline/regfile/data[23][29] ), .ip2(n18044), .s(
        n21596), .op(n9163) );
  mux2_1 U20140 ( .ip1(\pipeline/regfile/data[6][29] ), .ip2(n18044), .s(
        n21597), .op(n9707) );
  mux2_1 U20141 ( .ip1(\pipeline/regfile/data[5][29] ), .ip2(n18044), .s(
        n21598), .op(n9739) );
  mux2_1 U20142 ( .ip1(\pipeline/regfile/data[3][29] ), .ip2(n18044), .s(
        n21599), .op(n9803) );
  mux2_1 U20143 ( .ip1(\pipeline/regfile/data[13][29] ), .ip2(n18044), .s(
        n21600), .op(n9483) );
  mux2_1 U20144 ( .ip1(\pipeline/regfile/data[20][29] ), .ip2(n18044), .s(
        n21601), .op(n9259) );
  mux2_1 U20145 ( .ip1(\pipeline/regfile/data[25][29] ), .ip2(n18044), .s(
        n21602), .op(n9099) );
  mux2_1 U20146 ( .ip1(\pipeline/regfile/data[24][29] ), .ip2(n18044), .s(
        n21603), .op(n9131) );
  mux2_1 U20147 ( .ip1(\pipeline/regfile/data[14][29] ), .ip2(n18044), .s(
        n21604), .op(n9451) );
  mux2_1 U20148 ( .ip1(\pipeline/regfile/data[4][29] ), .ip2(n18044), .s(
        n21605), .op(n9771) );
  mux2_1 U20149 ( .ip1(\pipeline/regfile/data[31][29] ), .ip2(n18044), .s(
        n21606), .op(n8907) );
  mux2_1 U20150 ( .ip1(\pipeline/regfile/data[26][29] ), .ip2(n18044), .s(
        n21607), .op(n9067) );
  mux2_1 U20151 ( .ip1(\pipeline/regfile/data[16][29] ), .ip2(n18044), .s(
        n21608), .op(n9387) );
  mux2_1 U20152 ( .ip1(\pipeline/regfile/data[9][29] ), .ip2(n18044), .s(
        n21609), .op(n9611) );
  mux2_1 U20153 ( .ip1(\pipeline/regfile/data[2][29] ), .ip2(n18044), .s(
        n21610), .op(n9835) );
  mux2_1 U20154 ( .ip1(\pipeline/regfile/data[1][29] ), .ip2(n18044), .s(
        n21611), .op(n9867) );
  mux2_1 U20155 ( .ip1(\pipeline/regfile/data[27][29] ), .ip2(n18044), .s(
        n21612), .op(n9035) );
  mux2_1 U20156 ( .ip1(\pipeline/regfile/data[15][29] ), .ip2(n18044), .s(
        n21613), .op(n9419) );
  mux2_1 U20157 ( .ip1(\pipeline/regfile/data[7][29] ), .ip2(n18044), .s(
        n21614), .op(n9675) );
  mux2_1 U20158 ( .ip1(\pipeline/regfile/data[21][29] ), .ip2(n18044), .s(
        n21615), .op(n9227) );
  mux2_1 U20159 ( .ip1(\pipeline/regfile/data[17][29] ), .ip2(n18044), .s(
        n21616), .op(n9355) );
  mux2_1 U20160 ( .ip1(\pipeline/regfile/data[8][29] ), .ip2(n18044), .s(
        n21617), .op(n9643) );
  mux2_1 U20161 ( .ip1(\pipeline/regfile/data[10][29] ), .ip2(n18044), .s(
        n21618), .op(n9579) );
  mux2_1 U20162 ( .ip1(\pipeline/regfile/data[29][29] ), .ip2(n18044), .s(
        n21619), .op(n8971) );
  nand2_1 U20163 ( .ip1(\pipeline/csr/from_host [13]), .ip2(n22372), .op(
        n18046) );
  nand2_1 U20164 ( .ip1(n22373), .ip2(n22166), .op(n18045) );
  nand2_1 U20165 ( .ip1(n18046), .ip2(n18045), .op(n9947) );
  nand2_1 U20166 ( .ip1(n22378), .ip2(n22166), .op(n18048) );
  nand2_1 U20167 ( .ip1(\pipeline/csr/to_host [13]), .ip2(n22376), .op(n18047)
         );
  nand2_1 U20168 ( .ip1(n18048), .ip2(n18047), .op(n8759) );
  nand2_1 U20169 ( .ip1(\pipeline/csr/mtimecmp [13]), .ip2(n22363), .op(n18050) );
  nand2_1 U20170 ( .ip1(n22365), .ip2(n22166), .op(n18049) );
  nand2_1 U20171 ( .ip1(n18050), .ip2(n18049), .op(n10009) );
  inv_1 U20172 ( .ip(\pipeline/csr/instret_full [13]), .op(n18052) );
  nor2_1 U20173 ( .ip1(n18052), .ip2(n20990), .op(n18055) );
  mux2_1 U20174 ( .ip1(n18052), .ip2(\pipeline/csr/instret_full [13]), .s(
        n18051), .op(n18053) );
  nor2_1 U20175 ( .ip1(n21005), .ip2(n18053), .op(n18054) );
  ab_or_c_or_d U20176 ( .ip1(n21019), .ip2(n22166), .ip3(n18055), .ip4(n18054), 
        .op(n10125) );
  inv_1 U20177 ( .ip(n22166), .op(n20270) );
  nor2_1 U20178 ( .ip1(n20270), .ip2(n21168), .op(n18060) );
  inv_1 U20179 ( .ip(\pipeline/PC_WB [13]), .op(n18058) );
  inv_1 U20180 ( .ip(n20699), .op(n18056) );
  nand2_1 U20181 ( .ip1(n18056), .ip2(\pipeline/PC_WB [12]), .op(n18057) );
  not_ab_or_c_or_d U20182 ( .ip1(n18058), .ip2(n18057), .ip3(n19839), .ip4(
        n21171), .op(n18059) );
  ab_or_c_or_d U20183 ( .ip1(n21174), .ip2(\pipeline/epc [13]), .ip3(n18060), 
        .ip4(n18059), .op(n8858) );
  nand2_1 U20184 ( .ip1(n21032), .ip2(n22166), .op(n18062) );
  nand2_1 U20185 ( .ip1(\pipeline/csr/mtvec [13]), .ip2(n20705), .op(n18061)
         );
  nand2_1 U20186 ( .ip1(n18062), .ip2(n18061), .op(n9979) );
  nor2_1 U20187 ( .ip1(n18068), .ip2(n18067), .op(n18063) );
  nor2_1 U20188 ( .ip1(n18063), .ip2(n22665), .op(n18064) );
  nor2_1 U20189 ( .ip1(n18216), .ip2(n18064), .op(n18066) );
  nor2_1 U20190 ( .ip1(n18066), .ip2(n18065), .op(n18070) );
  nor4_1 U20191 ( .ip1(\pipeline/md_resp_result [11]), .ip2(n18068), .ip3(
        n18067), .ip4(n18219), .op(n18069) );
  not_ab_or_c_or_d U20192 ( .ip1(n18211), .ip2(n20554), .ip3(n18070), .ip4(
        n18069), .op(n18088) );
  not_ab_or_c_or_d U20193 ( .ip1(\pipeline/md/result [43]), .ip2(n18072), 
        .ip3(n18071), .ip4(n21505), .op(n18080) );
  or2_1 U20194 ( .ip1(n18073), .ip2(n18082), .op(n18078) );
  nand3_1 U20195 ( .ip1(n18075), .ip2(n18074), .ip3(n18081), .op(n18076) );
  or2_1 U20196 ( .ip1(n18076), .ip2(n18082), .op(n18077) );
  nand2_1 U20197 ( .ip1(n18078), .ip2(n18077), .op(n18079) );
  not_ab_or_c_or_d U20198 ( .ip1(\pipeline/md/result [43]), .ip2(n21509), 
        .ip3(n18080), .ip4(n18079), .op(n18085) );
  nand3_1 U20199 ( .ip1(n18083), .ip2(n18082), .ip3(n18081), .op(n18084) );
  nand2_1 U20200 ( .ip1(n18085), .ip2(n18084), .op(n18086) );
  nand2_1 U20201 ( .ip1(n20552), .ip2(n18086), .op(n18087) );
  nand2_1 U20202 ( .ip1(n18088), .ip2(n18087), .op(n18089) );
  mux2_1 U20203 ( .ip1(n18089), .ip2(\pipeline/md_resp_result [11]), .s(n21517), .op(n8623) );
  nand2_1 U20204 ( .ip1(n21032), .ip2(n22156), .op(n18091) );
  nand2_1 U20205 ( .ip1(\pipeline/csr/mtvec [11]), .ip2(n20705), .op(n18090)
         );
  nand2_1 U20206 ( .ip1(n18091), .ip2(n18090), .op(n9981) );
  nand2_1 U20207 ( .ip1(\pipeline/csr/from_host [11]), .ip2(n22372), .op(
        n18093) );
  nand2_1 U20208 ( .ip1(n22373), .ip2(n22156), .op(n18092) );
  nand2_1 U20209 ( .ip1(n18093), .ip2(n18092), .op(n9949) );
  nand2_1 U20210 ( .ip1(n22378), .ip2(n22156), .op(n18095) );
  nand2_1 U20211 ( .ip1(\pipeline/csr/to_host [11]), .ip2(n22376), .op(n18094)
         );
  nand2_1 U20212 ( .ip1(n18095), .ip2(n18094), .op(n8761) );
  nand2_1 U20213 ( .ip1(\pipeline/csr/mtimecmp [11]), .ip2(n22363), .op(n18097) );
  nand2_1 U20214 ( .ip1(n22365), .ip2(n22156), .op(n18096) );
  nand2_1 U20215 ( .ip1(n18097), .ip2(n18096), .op(n10011) );
  nor2_1 U20216 ( .ip1(n18838), .ip2(n18098), .op(n20461) );
  inv_1 U20217 ( .ip(n18110), .op(n18099) );
  nor4_1 U20218 ( .ip1(\pipeline/md_resp_result [22]), .ip2(n18109), .ip3(
        n18099), .ip4(n22755), .op(n18108) );
  not_ab_or_c_or_d U20219 ( .ip1(\pipeline/md/result [54]), .ip2(n18100), 
        .ip3(n18117), .ip4(n21505), .op(n18105) );
  nor2_1 U20220 ( .ip1(n18101), .ip2(n21659), .op(n18103) );
  nor2_1 U20221 ( .ip1(n18122), .ip2(n18103), .op(n18102) );
  not_ab_or_c_or_d U20222 ( .ip1(n18122), .ip2(n18103), .ip3(n21960), .ip4(
        n18102), .op(n18104) );
  not_ab_or_c_or_d U20223 ( .ip1(n21509), .ip2(\pipeline/md/result [54]), 
        .ip3(n18105), .ip4(n18104), .op(n18106) );
  nor2_1 U20224 ( .ip1(n18106), .ip2(n21967), .op(n18107) );
  not_ab_or_c_or_d U20225 ( .ip1(n20306), .ip2(n20461), .ip3(n18108), .ip4(
        n18107), .op(n18116) );
  inv_1 U20226 ( .ip(n18109), .op(n18111) );
  nand2_1 U20227 ( .ip1(n18111), .ip2(n18110), .op(n18112) );
  nand2_1 U20228 ( .ip1(n20310), .ip2(n18112), .op(n18113) );
  nand2_1 U20229 ( .ip1(n22738), .ip2(n18113), .op(n18114) );
  nand2_1 U20230 ( .ip1(\pipeline/md_resp_result [22]), .ip2(n18114), .op(
        n18115) );
  nand2_1 U20231 ( .ip1(n18116), .ip2(n18115), .op(n8612) );
  nor2_1 U20232 ( .ip1(n18117), .ip2(n21659), .op(n18119) );
  nor2_1 U20233 ( .ip1(\pipeline/md/result [55]), .ip2(n18119), .op(n18118) );
  not_ab_or_c_or_d U20234 ( .ip1(\pipeline/md/result [55]), .ip2(n18119), 
        .ip3(n21662), .ip4(n18118), .op(n18127) );
  inv_1 U20235 ( .ip(n18120), .op(n18125) );
  nor3_1 U20236 ( .ip1(n21957), .ip2(n18122), .ip3(n18121), .op(n18123) );
  nor3_1 U20237 ( .ip1(n20669), .ip2(n18125), .ip3(n18123), .op(n18124) );
  not_ab_or_c_or_d U20238 ( .ip1(n18125), .ip2(n21957), .ip3(n18124), .ip4(
        n21958), .op(n18126) );
  nor2_1 U20239 ( .ip1(n18127), .ip2(n18126), .op(n18128) );
  nor2_1 U20240 ( .ip1(n18128), .ip2(n21967), .op(n18130) );
  nor4_1 U20241 ( .ip1(\pipeline/md_resp_result [23]), .ip2(n18132), .ip3(
        n18131), .ip4(n22755), .op(n18129) );
  not_ab_or_c_or_d U20242 ( .ip1(n20461), .ip2(n21671), .ip3(n18130), .ip4(
        n18129), .op(n18137) );
  or2_1 U20243 ( .ip1(n18132), .ip2(n18131), .op(n18133) );
  nand2_1 U20244 ( .ip1(n20310), .ip2(n18133), .op(n18134) );
  nand2_1 U20245 ( .ip1(n22738), .ip2(n18134), .op(n18135) );
  nand2_1 U20246 ( .ip1(\pipeline/md_resp_result [23]), .ip2(n18135), .op(
        n18136) );
  nand2_1 U20247 ( .ip1(n18137), .ip2(n18136), .op(n8611) );
  nand2_1 U20248 ( .ip1(\pipeline/csr/from_host [17]), .ip2(n22372), .op(
        n18139) );
  nand2_1 U20249 ( .ip1(n22373), .ip2(n22183), .op(n18138) );
  nand2_1 U20250 ( .ip1(n18139), .ip2(n18138), .op(n9943) );
  nand2_1 U20251 ( .ip1(n22378), .ip2(n22183), .op(n18141) );
  nand2_1 U20252 ( .ip1(\pipeline/csr/to_host [17]), .ip2(n22376), .op(n18140)
         );
  nand2_1 U20253 ( .ip1(n18141), .ip2(n18140), .op(n8755) );
  nand2_1 U20254 ( .ip1(\pipeline/csr/mtimecmp [17]), .ip2(n22363), .op(n18143) );
  nand2_1 U20255 ( .ip1(n22365), .ip2(n22183), .op(n18142) );
  nand2_1 U20256 ( .ip1(n18143), .ip2(n18142), .op(n10005) );
  and3_1 U20257 ( .ip1(n20965), .ip2(n18144), .ip3(n20966), .op(n22357) );
  nor2_1 U20258 ( .ip1(htif_reset), .ip2(n22357), .op(n22356) );
  nand2_1 U20259 ( .ip1(\pipeline/csr/mie [17]), .ip2(n22356), .op(n18146) );
  nand2_1 U20260 ( .ip1(n22357), .ip2(n22183), .op(n18145) );
  nand2_1 U20261 ( .ip1(n18146), .ip2(n18145), .op(n10043) );
  inv_1 U20262 ( .ip(n20649), .op(n20633) );
  nor2_1 U20263 ( .ip1(n21499), .ip2(n20430), .op(n18147) );
  nor2_1 U20264 ( .ip1(n20633), .ip2(n18147), .op(n18150) );
  inv_1 U20265 ( .ip(n20647), .op(n20634) );
  nand2_1 U20266 ( .ip1(n20634), .ip2(n20430), .op(n18149) );
  mux2_1 U20267 ( .ip1(n18150), .ip2(n18149), .s(n18148), .op(n18156) );
  xor2_1 U20268 ( .ip1(\pipeline/md/b [16]), .ip2(n18151), .op(n18152) );
  nor2_1 U20269 ( .ip1(n21884), .ip2(n18152), .op(n18153) );
  xor2_1 U20270 ( .ip1(\pipeline/md/a [16]), .ip2(n18153), .op(n18154) );
  nand2_1 U20271 ( .ip1(n18154), .ip2(n21643), .op(n18155) );
  nand2_1 U20272 ( .ip1(n18156), .ip2(n18155), .op(n8425) );
  nand2_1 U20273 ( .ip1(\pipeline/md/negate_output ), .ip2(n18157), .op(n18158) );
  nand2_1 U20274 ( .ip1(n18159), .ip2(n18158), .op(n18161) );
  nor2_1 U20275 ( .ip1(n18162), .ip2(n18161), .op(n18160) );
  not_ab_or_c_or_d U20276 ( .ip1(n18162), .ip2(n18161), .ip3(n21960), .ip4(
        n18160), .op(n18169) );
  nor2_1 U20277 ( .ip1(\pipeline/md/result [45]), .ip2(n18163), .op(n18164) );
  nor3_1 U20278 ( .ip1(\pipeline/md/result [46]), .ip2(n18164), .ip3(n21966), 
        .op(n18167) );
  inv_1 U20279 ( .ip(n18164), .op(n18165) );
  inv_1 U20280 ( .ip(\pipeline/md/result [46]), .op(n22611) );
  not_ab_or_c_or_d U20281 ( .ip1(\pipeline/md/negate_output ), .ip2(n18165), 
        .ip3(n22611), .ip4(n21967), .op(n18166) );
  nor3_1 U20282 ( .ip1(n21972), .ip2(n18167), .ip3(n18166), .op(n18168) );
  nor2_1 U20283 ( .ip1(n18169), .ip2(n18168), .op(n18173) );
  nor3_1 U20284 ( .ip1(n18171), .ip2(n22755), .ip3(n18170), .op(n18172) );
  not_ab_or_c_or_d U20285 ( .ip1(n20306), .ip2(n18174), .ip3(n18173), .ip4(
        n18172), .op(n18181) );
  nand2_1 U20286 ( .ip1(n18176), .ip2(n18175), .op(n18177) );
  nand2_1 U20287 ( .ip1(n20310), .ip2(n18177), .op(n18178) );
  nand2_1 U20288 ( .ip1(n22738), .ip2(n18178), .op(n18179) );
  nand2_1 U20289 ( .ip1(\pipeline/md_resp_result [14]), .ip2(n18179), .op(
        n18180) );
  nand2_1 U20290 ( .ip1(n18181), .ip2(n18180), .op(n8620) );
  nor2_1 U20291 ( .ip1(n18182), .ip2(n21659), .op(n18183) );
  xor2_1 U20292 ( .ip1(n18184), .ip2(n18183), .op(n18185) );
  nor2_1 U20293 ( .ip1(n21960), .ip2(n18185), .op(n18189) );
  not_ab_or_c_or_d U20294 ( .ip1(\pipeline/md/result [48]), .ip2(n18187), 
        .ip3(n21662), .ip4(n18186), .op(n18188) );
  not_ab_or_c_or_d U20295 ( .ip1(n21509), .ip2(\pipeline/md/result [48]), 
        .ip3(n18189), .ip4(n18188), .op(n18190) );
  nor2_1 U20296 ( .ip1(n18190), .ip2(n21967), .op(n18200) );
  nor2_1 U20297 ( .ip1(n18196), .ip2(n18195), .op(n18191) );
  nor2_1 U20298 ( .ip1(n18191), .ip2(n22665), .op(n18192) );
  nor2_1 U20299 ( .ip1(n18216), .ip2(n18192), .op(n18194) );
  nor2_1 U20300 ( .ip1(n18194), .ip2(n18193), .op(n18199) );
  nor4_1 U20301 ( .ip1(\pipeline/md_resp_result [16]), .ip2(n18196), .ip3(
        n18195), .ip4(n18219), .op(n18198) );
  nor2_1 U20302 ( .ip1(n21516), .ip2(n18838), .op(n18197) );
  or4_1 U20303 ( .ip1(n18200), .ip2(n18199), .ip3(n18198), .ip4(n18197), .op(
        n18201) );
  mux2_1 U20304 ( .ip1(n18201), .ip2(\pipeline/md_resp_result [16]), .s(n21517), .op(n8618) );
  nor2_1 U20305 ( .ip1(n18202), .ip2(n21659), .op(n18203) );
  mux2_1 U20306 ( .ip1(n18204), .ip2(\pipeline/md/result [40]), .s(n18203), 
        .op(n18210) );
  nor2_1 U20307 ( .ip1(n18205), .ip2(n21659), .op(n18207) );
  nor2_1 U20308 ( .ip1(n18208), .ip2(n18207), .op(n18206) );
  not_ab_or_c_or_d U20309 ( .ip1(n18208), .ip2(n18207), .ip3(n21960), .ip4(
        n18206), .op(n18209) );
  not_ab_or_c_or_d U20310 ( .ip1(n21960), .ip2(n18210), .ip3(n18209), .ip4(
        n21967), .op(n18225) );
  inv_1 U20311 ( .ip(n18211), .op(n18212) );
  nor2_1 U20312 ( .ip1(n18213), .ip2(n18212), .op(n18224) );
  nor2_1 U20313 ( .ip1(n18221), .ip2(n18220), .op(n18214) );
  nor2_1 U20314 ( .ip1(n18214), .ip2(n22665), .op(n18215) );
  nor2_1 U20315 ( .ip1(n18216), .ip2(n18215), .op(n18218) );
  nor2_1 U20316 ( .ip1(n18218), .ip2(n18217), .op(n18223) );
  nor4_1 U20317 ( .ip1(\pipeline/md_resp_result [8]), .ip2(n18221), .ip3(
        n18220), .ip4(n18219), .op(n18222) );
  or4_1 U20318 ( .ip1(n18225), .ip2(n18224), .ip3(n18223), .ip4(n18222), .op(
        n18226) );
  mux2_1 U20319 ( .ip1(n18226), .ip2(\pipeline/md_resp_result [8]), .s(n21517), 
        .op(n8626) );
  nand2_1 U20320 ( .ip1(n18228), .ip2(n18227), .op(n18236) );
  inv_1 U20321 ( .ip(n18229), .op(n18230) );
  nand2_1 U20322 ( .ip1(n18231), .ip2(n18230), .op(n18234) );
  inv_1 U20323 ( .ip(n18232), .op(n18233) );
  nand2_1 U20324 ( .ip1(n18234), .ip2(n18233), .op(n18235) );
  xnor2_1 U20325 ( .ip1(n18236), .ip2(n18235), .op(imem_haddr[7]) );
  nand2_1 U20326 ( .ip1(n21995), .ip2(imem_haddr[7]), .op(n18238) );
  nand2_1 U20327 ( .ip1(\pipeline/PC_IF [7]), .ip2(n21996), .op(n18237) );
  nand2_1 U20328 ( .ip1(n18238), .ip2(n18237), .op(n8476) );
  nand2_1 U20329 ( .ip1(\pipeline/PC_IF [7]), .ip2(n22048), .op(n18240) );
  nand2_1 U20330 ( .ip1(\pipeline/PC_DX [7]), .ip2(n21999), .op(n18239) );
  nand2_1 U20331 ( .ip1(n18240), .ip2(n18239), .op(n8475) );
  mux2_1 U20332 ( .ip1(\pipeline/PC_WB [7]), .ip2(\pipeline/PC_DX [7]), .s(
        n22067), .op(n8896) );
  nand2_1 U20333 ( .ip1(n21032), .ip2(n19677), .op(n18242) );
  nand2_1 U20334 ( .ip1(\pipeline/csr/mtvec [7]), .ip2(n20705), .op(n18241) );
  nand2_1 U20335 ( .ip1(n18242), .ip2(n18241), .op(n9985) );
  nand2_1 U20336 ( .ip1(n18243), .ip2(n21583), .op(n18244) );
  nand2_1 U20337 ( .ip1(n18245), .ip2(n18244), .op(n18246) );
  buf_1 U20338 ( .ip(n21619), .op(n19353) );
  mux2_1 U20339 ( .ip1(\pipeline/regfile/data[29][7] ), .ip2(n18246), .s(
        n19353), .op(n8993) );
  buf_1 U20340 ( .ip(n21604), .op(n19354) );
  mux2_1 U20341 ( .ip1(\pipeline/regfile/data[14][7] ), .ip2(n18246), .s(
        n19354), .op(n9473) );
  buf_1 U20342 ( .ip(n21589), .op(n19355) );
  mux2_1 U20343 ( .ip1(\pipeline/regfile/data[22][7] ), .ip2(n18246), .s(
        n19355), .op(n9217) );
  buf_1 U20344 ( .ip(n21598), .op(n19356) );
  mux2_1 U20345 ( .ip1(\pipeline/regfile/data[5][7] ), .ip2(n18246), .s(n19356), .op(n9761) );
  buf_1 U20346 ( .ip(n21612), .op(n19357) );
  mux2_1 U20347 ( .ip1(\pipeline/regfile/data[27][7] ), .ip2(n18246), .s(
        n19357), .op(n9057) );
  buf_1 U20348 ( .ip(n21607), .op(n19358) );
  mux2_1 U20349 ( .ip1(\pipeline/regfile/data[26][7] ), .ip2(n18246), .s(
        n19358), .op(n9089) );
  buf_1 U20350 ( .ip(n21590), .op(n19359) );
  mux2_1 U20351 ( .ip1(\pipeline/regfile/data[28][7] ), .ip2(n18246), .s(
        n19359), .op(n9025) );
  buf_1 U20352 ( .ip(n21606), .op(n19360) );
  mux2_1 U20353 ( .ip1(\pipeline/regfile/data[31][7] ), .ip2(n18246), .s(
        n19360), .op(n8929) );
  buf_1 U20354 ( .ip(n21592), .op(n19361) );
  mux2_1 U20355 ( .ip1(\pipeline/regfile/data[19][7] ), .ip2(n18246), .s(
        n19361), .op(n9313) );
  buf_1 U20356 ( .ip(n21597), .op(n19362) );
  mux2_1 U20357 ( .ip1(\pipeline/regfile/data[6][7] ), .ip2(n18246), .s(n19362), .op(n9729) );
  buf_1 U20358 ( .ip(n21594), .op(n19363) );
  mux2_1 U20359 ( .ip1(\pipeline/regfile/data[30][7] ), .ip2(n18246), .s(
        n19363), .op(n8961) );
  buf_1 U20360 ( .ip(n21595), .op(n19364) );
  mux2_1 U20361 ( .ip1(\pipeline/regfile/data[18][7] ), .ip2(n18246), .s(
        n19364), .op(n9345) );
  buf_1 U20362 ( .ip(n21593), .op(n19365) );
  mux2_1 U20363 ( .ip1(\pipeline/regfile/data[11][7] ), .ip2(n18246), .s(
        n19365), .op(n9569) );
  buf_1 U20364 ( .ip(n21602), .op(n19366) );
  mux2_1 U20365 ( .ip1(\pipeline/regfile/data[25][7] ), .ip2(n18246), .s(
        n19366), .op(n9121) );
  buf_1 U20366 ( .ip(n21600), .op(n19367) );
  mux2_1 U20367 ( .ip1(\pipeline/regfile/data[13][7] ), .ip2(n18246), .s(
        n19367), .op(n9505) );
  buf_1 U20368 ( .ip(n21616), .op(n19368) );
  mux2_1 U20369 ( .ip1(\pipeline/regfile/data[17][7] ), .ip2(n18246), .s(
        n19368), .op(n9377) );
  buf_1 U20370 ( .ip(n21596), .op(n19369) );
  mux2_1 U20371 ( .ip1(\pipeline/regfile/data[23][7] ), .ip2(n18246), .s(
        n19369), .op(n9185) );
  buf_1 U20372 ( .ip(n21591), .op(n19370) );
  mux2_1 U20373 ( .ip1(\pipeline/regfile/data[12][7] ), .ip2(n18246), .s(
        n19370), .op(n9537) );
  buf_1 U20374 ( .ip(n21614), .op(n19371) );
  mux2_1 U20375 ( .ip1(\pipeline/regfile/data[7][7] ), .ip2(n18246), .s(n19371), .op(n9697) );
  buf_1 U20376 ( .ip(n21617), .op(n19372) );
  mux2_1 U20377 ( .ip1(\pipeline/regfile/data[8][7] ), .ip2(n18246), .s(n19372), .op(n9665) );
  buf_1 U20378 ( .ip(n21613), .op(n19373) );
  mux2_1 U20379 ( .ip1(\pipeline/regfile/data[15][7] ), .ip2(n18246), .s(
        n19373), .op(n9441) );
  buf_1 U20380 ( .ip(n21618), .op(n19374) );
  mux2_1 U20381 ( .ip1(\pipeline/regfile/data[10][7] ), .ip2(n18246), .s(
        n19374), .op(n9601) );
  buf_1 U20382 ( .ip(n21615), .op(n19375) );
  mux2_1 U20383 ( .ip1(\pipeline/regfile/data[21][7] ), .ip2(n18246), .s(
        n19375), .op(n9249) );
  buf_1 U20384 ( .ip(n21603), .op(n19376) );
  mux2_1 U20385 ( .ip1(\pipeline/regfile/data[24][7] ), .ip2(n18246), .s(
        n19376), .op(n9153) );
  buf_1 U20386 ( .ip(n21601), .op(n19377) );
  mux2_1 U20387 ( .ip1(\pipeline/regfile/data[20][7] ), .ip2(n18246), .s(
        n19377), .op(n9281) );
  buf_1 U20388 ( .ip(n21609), .op(n19378) );
  mux2_1 U20389 ( .ip1(\pipeline/regfile/data[9][7] ), .ip2(n18246), .s(n19378), .op(n9633) );
  buf_1 U20390 ( .ip(n21608), .op(n19379) );
  mux2_1 U20391 ( .ip1(\pipeline/regfile/data[16][7] ), .ip2(n18246), .s(
        n19379), .op(n9409) );
  buf_1 U20392 ( .ip(n21599), .op(n19380) );
  mux2_1 U20393 ( .ip1(\pipeline/regfile/data[3][7] ), .ip2(n18246), .s(n19380), .op(n9825) );
  buf_1 U20394 ( .ip(n21611), .op(n19381) );
  mux2_1 U20395 ( .ip1(\pipeline/regfile/data[1][7] ), .ip2(n18246), .s(n19381), .op(n9889) );
  buf_1 U20396 ( .ip(n21610), .op(n19382) );
  mux2_1 U20397 ( .ip1(\pipeline/regfile/data[2][7] ), .ip2(n18246), .s(n19382), .op(n9857) );
  buf_1 U20398 ( .ip(n21605), .op(n19383) );
  mux2_1 U20399 ( .ip1(\pipeline/regfile/data[4][7] ), .ip2(n18246), .s(n19383), .op(n9793) );
  nor2_1 U20400 ( .ip1(n22274), .ip2(n21029), .op(n18250) );
  inv_1 U20401 ( .ip(\pipeline/csr/mtvec [23]), .op(n18247) );
  nor2_1 U20402 ( .ip1(htif_reset), .ip2(n18247), .op(n18248) );
  nor2_1 U20403 ( .ip1(n21032), .ip2(n18248), .op(n18249) );
  nor2_1 U20404 ( .ip1(n18250), .ip2(n18249), .op(n9969) );
  nor4_1 U20405 ( .ip1(\pipeline/md_resp_result [20]), .ip2(n18263), .ip3(
        n18264), .ip4(n22755), .op(n18262) );
  nor2_1 U20406 ( .ip1(n18251), .ip2(n21659), .op(n18254) );
  nor2_1 U20407 ( .ip1(n18253), .ip2(n18254), .op(n18252) );
  not_ab_or_c_or_d U20408 ( .ip1(n18254), .ip2(n18253), .ip3(n21960), .ip4(
        n18252), .op(n18260) );
  inv_1 U20409 ( .ip(n18256), .op(n18255) );
  nor3_1 U20410 ( .ip1(\pipeline/md/result [52]), .ip2(n21966), .ip3(n18255), 
        .op(n18258) );
  inv_1 U20411 ( .ip(\pipeline/md/result [52]), .op(n22669) );
  not_ab_or_c_or_d U20412 ( .ip1(\pipeline/md/negate_output ), .ip2(n18256), 
        .ip3(n22669), .ip4(n21967), .op(n18257) );
  nor3_1 U20413 ( .ip1(n21972), .ip2(n18258), .ip3(n18257), .op(n18259) );
  nor2_1 U20414 ( .ip1(n18260), .ip2(n18259), .op(n18261) );
  not_ab_or_c_or_d U20415 ( .ip1(n20461), .ip2(n21977), .ip3(n18262), .ip4(
        n18261), .op(n18269) );
  or2_1 U20416 ( .ip1(n18264), .ip2(n18263), .op(n18265) );
  nand2_1 U20417 ( .ip1(n20310), .ip2(n18265), .op(n18266) );
  nand2_1 U20418 ( .ip1(n22738), .ip2(n18266), .op(n18267) );
  nand2_1 U20419 ( .ip1(\pipeline/md_resp_result [20]), .ip2(n18267), .op(
        n18268) );
  nand2_1 U20420 ( .ip1(n18269), .ip2(n18268), .op(n8614) );
  nand2_1 U20421 ( .ip1(n21032), .ip2(n22183), .op(n18271) );
  nand2_1 U20422 ( .ip1(\pipeline/csr/mtvec [17]), .ip2(n20705), .op(n18270)
         );
  nand2_1 U20423 ( .ip1(n18271), .ip2(n18270), .op(n9975) );
  nand2_1 U20424 ( .ip1(n21043), .ip2(n22177), .op(n18276) );
  inv_1 U20425 ( .ip(n18272), .op(n19902) );
  xor2_1 U20426 ( .ip1(n19902), .ip2(\pipeline/PC_WB [15]), .op(n18273) );
  nand2_1 U20427 ( .ip1(n21046), .ip2(n18273), .op(n18275) );
  nand2_1 U20428 ( .ip1(\pipeline/epc [15]), .ip2(n21174), .op(n18274) );
  nand3_1 U20429 ( .ip1(n18276), .ip2(n18275), .ip3(n18274), .op(n8856) );
  nor2_1 U20430 ( .ip1(n21029), .ip2(n22177), .op(n18280) );
  inv_1 U20431 ( .ip(\pipeline/csr/mtvec [15]), .op(n18277) );
  nor2_1 U20432 ( .ip1(htif_reset), .ip2(n18277), .op(n18278) );
  nor2_1 U20433 ( .ip1(n21032), .ip2(n18278), .op(n18279) );
  nor2_1 U20434 ( .ip1(n18280), .ip2(n18279), .op(n9977) );
  mux2_1 U20435 ( .ip1(\pipeline/dmem_type_WB [0]), .ip2(dmem_hsize[0]), .s(
        n19498), .op(n8775) );
  nor2_1 U20436 ( .ip1(\pipeline/dmem_type_WB [1]), .ip2(
        \pipeline/dmem_type_WB [0]), .op(n22071) );
  nor3_1 U20437 ( .ip1(n22071), .ip2(n18281), .ip3(n21583), .op(n18282) );
  ab_or_c_or_d U20438 ( .ip1(n18283), .ip2(n21583), .ip3(n18282), .ip4(n19390), 
        .op(n18284) );
  mux2_1 U20439 ( .ip1(\pipeline/regfile/data[29][15] ), .ip2(n18284), .s(
        n21619), .op(n8985) );
  mux2_1 U20440 ( .ip1(\pipeline/regfile/data[14][15] ), .ip2(n18284), .s(
        n21604), .op(n9465) );
  mux2_1 U20441 ( .ip1(\pipeline/regfile/data[22][15] ), .ip2(n18284), .s(
        n21589), .op(n9209) );
  mux2_1 U20442 ( .ip1(\pipeline/regfile/data[5][15] ), .ip2(n18284), .s(
        n21598), .op(n9753) );
  mux2_1 U20443 ( .ip1(\pipeline/regfile/data[27][15] ), .ip2(n18284), .s(
        n21612), .op(n9049) );
  mux2_1 U20444 ( .ip1(\pipeline/regfile/data[26][15] ), .ip2(n18284), .s(
        n21607), .op(n9081) );
  mux2_1 U20445 ( .ip1(\pipeline/regfile/data[28][15] ), .ip2(n18284), .s(
        n21590), .op(n9017) );
  mux2_1 U20446 ( .ip1(\pipeline/regfile/data[31][15] ), .ip2(n18284), .s(
        n21606), .op(n8921) );
  mux2_1 U20447 ( .ip1(\pipeline/regfile/data[19][15] ), .ip2(n18284), .s(
        n21592), .op(n9305) );
  mux2_1 U20448 ( .ip1(\pipeline/regfile/data[6][15] ), .ip2(n18284), .s(
        n21597), .op(n9721) );
  mux2_1 U20449 ( .ip1(\pipeline/regfile/data[30][15] ), .ip2(n18284), .s(
        n21594), .op(n8953) );
  mux2_1 U20450 ( .ip1(\pipeline/regfile/data[18][15] ), .ip2(n18284), .s(
        n21595), .op(n9337) );
  mux2_1 U20451 ( .ip1(\pipeline/regfile/data[11][15] ), .ip2(n18284), .s(
        n21593), .op(n9561) );
  mux2_1 U20452 ( .ip1(\pipeline/regfile/data[25][15] ), .ip2(n18284), .s(
        n21602), .op(n9113) );
  mux2_1 U20453 ( .ip1(\pipeline/regfile/data[13][15] ), .ip2(n18284), .s(
        n21600), .op(n9497) );
  mux2_1 U20454 ( .ip1(\pipeline/regfile/data[17][15] ), .ip2(n18284), .s(
        n21616), .op(n9369) );
  mux2_1 U20455 ( .ip1(\pipeline/regfile/data[23][15] ), .ip2(n18284), .s(
        n21596), .op(n9177) );
  mux2_1 U20456 ( .ip1(\pipeline/regfile/data[12][15] ), .ip2(n18284), .s(
        n21591), .op(n9529) );
  mux2_1 U20457 ( .ip1(\pipeline/regfile/data[7][15] ), .ip2(n18284), .s(
        n21614), .op(n9689) );
  mux2_1 U20458 ( .ip1(\pipeline/regfile/data[8][15] ), .ip2(n18284), .s(
        n21617), .op(n9657) );
  mux2_1 U20459 ( .ip1(\pipeline/regfile/data[15][15] ), .ip2(n18284), .s(
        n21613), .op(n9433) );
  mux2_1 U20460 ( .ip1(\pipeline/regfile/data[10][15] ), .ip2(n18284), .s(
        n21618), .op(n9593) );
  mux2_1 U20461 ( .ip1(\pipeline/regfile/data[21][15] ), .ip2(n18284), .s(
        n21615), .op(n9241) );
  mux2_1 U20462 ( .ip1(\pipeline/regfile/data[24][15] ), .ip2(n18284), .s(
        n21603), .op(n9145) );
  mux2_1 U20463 ( .ip1(\pipeline/regfile/data[20][15] ), .ip2(n18284), .s(
        n21601), .op(n9273) );
  mux2_1 U20464 ( .ip1(\pipeline/regfile/data[9][15] ), .ip2(n18284), .s(
        n21609), .op(n9625) );
  mux2_1 U20465 ( .ip1(\pipeline/regfile/data[16][15] ), .ip2(n18284), .s(
        n21608), .op(n9401) );
  mux2_1 U20466 ( .ip1(\pipeline/regfile/data[3][15] ), .ip2(n18284), .s(
        n21599), .op(n9817) );
  mux2_1 U20467 ( .ip1(\pipeline/regfile/data[1][15] ), .ip2(n18284), .s(
        n21611), .op(n9881) );
  mux2_1 U20468 ( .ip1(\pipeline/regfile/data[2][15] ), .ip2(n18284), .s(
        n21610), .op(n9849) );
  mux2_1 U20469 ( .ip1(\pipeline/regfile/data[4][15] ), .ip2(n18284), .s(
        n21605), .op(n9785) );
  inv_1 U20470 ( .ip(n18285), .op(n18286) );
  nor2_1 U20471 ( .ip1(n18287), .ip2(n18286), .op(n18289) );
  xor2_1 U20472 ( .ip1(n18289), .ip2(n18288), .op(imem_haddr[16]) );
  nand2_1 U20473 ( .ip1(n21995), .ip2(imem_haddr[16]), .op(n18291) );
  nand2_1 U20474 ( .ip1(\pipeline/PC_IF [16]), .ip2(n21996), .op(n18290) );
  nand2_1 U20475 ( .ip1(n18291), .ip2(n18290), .op(n8458) );
  nand2_1 U20476 ( .ip1(\pipeline/PC_IF [16]), .ip2(n22048), .op(n18293) );
  nand2_1 U20477 ( .ip1(\pipeline/PC_DX [16]), .ip2(n21999), .op(n18292) );
  nand2_1 U20478 ( .ip1(n18293), .ip2(n18292), .op(n8457) );
  nand2_1 U20479 ( .ip1(n18295), .ip2(n18294), .op(n18304) );
  nand2_1 U20480 ( .ip1(n18297), .ip2(n18296), .op(n18298) );
  inv_1 U20481 ( .ip(n18298), .op(n18300) );
  nand2_2 U20482 ( .ip1(n18300), .ip2(n18299), .op(n20042) );
  nand2_1 U20483 ( .ip1(n20042), .ip2(n20019), .op(n18302) );
  inv_1 U20484 ( .ip(n20021), .op(n18301) );
  nand2_1 U20485 ( .ip1(n18302), .ip2(n18301), .op(n18303) );
  xnor2_1 U20486 ( .ip1(n18304), .ip2(n18303), .op(imem_haddr[19]) );
  nand2_1 U20487 ( .ip1(n21995), .ip2(imem_haddr[19]), .op(n18306) );
  nand2_1 U20488 ( .ip1(\pipeline/PC_IF [19]), .ip2(n21996), .op(n18305) );
  nand2_1 U20489 ( .ip1(n18306), .ip2(n18305), .op(n8452) );
  nand2_1 U20490 ( .ip1(\pipeline/PC_IF [19]), .ip2(n21988), .op(n18308) );
  nand2_1 U20491 ( .ip1(\pipeline/PC_DX [19]), .ip2(n21999), .op(n18307) );
  nand2_1 U20492 ( .ip1(n18308), .ip2(n18307), .op(n8451) );
  or2_1 U20493 ( .ip1(n20692), .ip2(n18309), .op(n18311) );
  xor2_1 U20494 ( .ip1(n18311), .ip2(n18310), .op(imem_haddr[10]) );
  nand2_1 U20495 ( .ip1(n21995), .ip2(imem_haddr[10]), .op(n18313) );
  nand2_1 U20496 ( .ip1(\pipeline/PC_IF [10]), .ip2(n21996), .op(n18312) );
  nand2_1 U20497 ( .ip1(n18313), .ip2(n18312), .op(n8470) );
  nand2_1 U20498 ( .ip1(\pipeline/PC_IF [10]), .ip2(n22048), .op(n18315) );
  nand2_1 U20499 ( .ip1(\pipeline/PC_DX [10]), .ip2(n21999), .op(n18314) );
  nand2_1 U20500 ( .ip1(n18315), .ip2(n18314), .op(n8469) );
  mux2_1 U20501 ( .ip1(\pipeline/PC_WB [24]), .ip2(\pipeline/PC_DX [24]), .s(
        n22067), .op(n8879) );
  nand2_1 U20502 ( .ip1(n21995), .ip2(imem_haddr[25]), .op(n18317) );
  nand2_1 U20503 ( .ip1(\pipeline/PC_IF [25]), .ip2(n21996), .op(n18316) );
  nand2_1 U20504 ( .ip1(n18317), .ip2(n18316), .op(n8440) );
  nand2_1 U20505 ( .ip1(\pipeline/PC_IF [25]), .ip2(n22048), .op(n18319) );
  nand2_1 U20506 ( .ip1(\pipeline/PC_DX [25]), .ip2(n21999), .op(n18318) );
  nand2_1 U20507 ( .ip1(n18319), .ip2(n18318), .op(n8439) );
  mux2_1 U20508 ( .ip1(\pipeline/PC_WB [25]), .ip2(\pipeline/PC_DX [25]), .s(
        n19498), .op(n8878) );
  nand2_1 U20509 ( .ip1(\pipeline/csr/from_host [25]), .ip2(n22372), .op(
        n18321) );
  nand2_1 U20510 ( .ip1(n22373), .ip2(n22217), .op(n18320) );
  nand2_1 U20511 ( .ip1(n18321), .ip2(n18320), .op(n9935) );
  nand2_1 U20512 ( .ip1(n22378), .ip2(n22217), .op(n18323) );
  nand2_1 U20513 ( .ip1(\pipeline/csr/to_host [25]), .ip2(n22376), .op(n18322)
         );
  nand2_1 U20514 ( .ip1(n18323), .ip2(n18322), .op(n8747) );
  nand2_1 U20515 ( .ip1(\pipeline/csr/mtimecmp [25]), .ip2(n22363), .op(n18325) );
  nand2_1 U20516 ( .ip1(n22365), .ip2(n22217), .op(n18324) );
  nand2_1 U20517 ( .ip1(n18325), .ip2(n18324), .op(n9997) );
  nand2_1 U20518 ( .ip1(\pipeline/csr/mie [25]), .ip2(n22356), .op(n18327) );
  nand2_1 U20519 ( .ip1(n22357), .ip2(n22217), .op(n18326) );
  nand2_1 U20520 ( .ip1(n18327), .ip2(n18326), .op(n10035) );
  nand2_1 U20521 ( .ip1(n18568), .ip2(n18328), .op(n22252) );
  inv_1 U20522 ( .ip(n22252), .op(n21177) );
  inv_1 U20523 ( .ip(n18757), .op(n18329) );
  nor2_1 U20524 ( .ip1(\pipeline/csr/time_full [25]), .ip2(n18329), .op(n18331) );
  nor3_1 U20525 ( .ip1(n21177), .ip2(n19097), .ip3(n18331), .op(n18330) );
  not_ab_or_c_or_d U20526 ( .ip1(n21179), .ip2(n22217), .ip3(n21217), .ip4(
        n18330), .op(n18334) );
  inv_1 U20527 ( .ip(n21210), .op(n21198) );
  nor2_1 U20528 ( .ip1(n18331), .ip2(n19097), .op(n18332) );
  nor2_1 U20529 ( .ip1(n21198), .ip2(n18332), .op(n18333) );
  nor2_1 U20530 ( .ip1(n18334), .ip2(n18333), .op(\pipeline/csr/N1962 ) );
  nand2_1 U20531 ( .ip1(\pipeline/csr/mscratch [25]), .ip2(n22013), .op(n18336) );
  nand2_1 U20532 ( .ip1(n22014), .ip2(n22217), .op(n18335) );
  nand2_1 U20533 ( .ip1(n18336), .ip2(n18335), .op(n9903) );
  nor2_1 U20534 ( .ip1(n22217), .ip2(n21029), .op(n18340) );
  inv_1 U20535 ( .ip(\pipeline/csr/mtvec [25]), .op(n18337) );
  nor2_1 U20536 ( .ip1(n21089), .ip2(n18337), .op(n18338) );
  nor2_1 U20537 ( .ip1(n21032), .ip2(n18338), .op(n18339) );
  nor2_1 U20538 ( .ip1(n18340), .ip2(n18339), .op(n9967) );
  nand2_1 U20539 ( .ip1(n18341), .ip2(n21583), .op(n18343) );
  nand2_1 U20540 ( .ip1(dmem_rdata[25]), .ip2(n21585), .op(n18342) );
  nand3_1 U20541 ( .ip1(n21588), .ip2(n18343), .ip3(n18342), .op(n18344) );
  mux2_1 U20542 ( .ip1(\pipeline/regfile/data[29][25] ), .ip2(n18344), .s(
        n19353), .op(n8975) );
  mux2_1 U20543 ( .ip1(\pipeline/regfile/data[14][25] ), .ip2(n18344), .s(
        n19354), .op(n9455) );
  mux2_1 U20544 ( .ip1(\pipeline/regfile/data[22][25] ), .ip2(n18344), .s(
        n19355), .op(n9199) );
  mux2_1 U20545 ( .ip1(\pipeline/regfile/data[5][25] ), .ip2(n18344), .s(
        n19356), .op(n9743) );
  mux2_1 U20546 ( .ip1(\pipeline/regfile/data[27][25] ), .ip2(n18344), .s(
        n19357), .op(n9039) );
  mux2_1 U20547 ( .ip1(\pipeline/regfile/data[26][25] ), .ip2(n18344), .s(
        n19358), .op(n9071) );
  mux2_1 U20548 ( .ip1(\pipeline/regfile/data[28][25] ), .ip2(n18344), .s(
        n19359), .op(n9007) );
  mux2_1 U20549 ( .ip1(\pipeline/regfile/data[31][25] ), .ip2(n18344), .s(
        n19360), .op(n8911) );
  mux2_1 U20550 ( .ip1(\pipeline/regfile/data[19][25] ), .ip2(n18344), .s(
        n19361), .op(n9295) );
  mux2_1 U20551 ( .ip1(\pipeline/regfile/data[6][25] ), .ip2(n18344), .s(
        n19362), .op(n9711) );
  mux2_1 U20552 ( .ip1(\pipeline/regfile/data[30][25] ), .ip2(n18344), .s(
        n19363), .op(n8943) );
  mux2_1 U20553 ( .ip1(\pipeline/regfile/data[18][25] ), .ip2(n18344), .s(
        n19364), .op(n9327) );
  mux2_1 U20554 ( .ip1(\pipeline/regfile/data[11][25] ), .ip2(n18344), .s(
        n19365), .op(n9551) );
  mux2_1 U20555 ( .ip1(\pipeline/regfile/data[25][25] ), .ip2(n18344), .s(
        n19366), .op(n9103) );
  mux2_1 U20556 ( .ip1(\pipeline/regfile/data[13][25] ), .ip2(n18344), .s(
        n19367), .op(n9487) );
  mux2_1 U20557 ( .ip1(\pipeline/regfile/data[17][25] ), .ip2(n18344), .s(
        n19368), .op(n9359) );
  mux2_1 U20558 ( .ip1(\pipeline/regfile/data[23][25] ), .ip2(n18344), .s(
        n19369), .op(n9167) );
  mux2_1 U20559 ( .ip1(\pipeline/regfile/data[12][25] ), .ip2(n18344), .s(
        n19370), .op(n9519) );
  mux2_1 U20560 ( .ip1(\pipeline/regfile/data[7][25] ), .ip2(n18344), .s(
        n19371), .op(n9679) );
  mux2_1 U20561 ( .ip1(\pipeline/regfile/data[8][25] ), .ip2(n18344), .s(
        n19372), .op(n9647) );
  mux2_1 U20562 ( .ip1(\pipeline/regfile/data[15][25] ), .ip2(n18344), .s(
        n19373), .op(n9423) );
  mux2_1 U20563 ( .ip1(\pipeline/regfile/data[10][25] ), .ip2(n18344), .s(
        n19374), .op(n9583) );
  mux2_1 U20564 ( .ip1(\pipeline/regfile/data[21][25] ), .ip2(n18344), .s(
        n19375), .op(n9231) );
  mux2_1 U20565 ( .ip1(\pipeline/regfile/data[24][25] ), .ip2(n18344), .s(
        n19376), .op(n9135) );
  mux2_1 U20566 ( .ip1(\pipeline/regfile/data[20][25] ), .ip2(n18344), .s(
        n19377), .op(n9263) );
  mux2_1 U20567 ( .ip1(\pipeline/regfile/data[9][25] ), .ip2(n18344), .s(
        n19378), .op(n9615) );
  mux2_1 U20568 ( .ip1(\pipeline/regfile/data[16][25] ), .ip2(n18344), .s(
        n19379), .op(n9391) );
  mux2_1 U20569 ( .ip1(\pipeline/regfile/data[3][25] ), .ip2(n18344), .s(
        n19380), .op(n9807) );
  mux2_1 U20570 ( .ip1(\pipeline/regfile/data[1][25] ), .ip2(n18344), .s(
        n19381), .op(n9871) );
  mux2_1 U20571 ( .ip1(\pipeline/regfile/data[2][25] ), .ip2(n18344), .s(
        n19382), .op(n9839) );
  mux2_1 U20572 ( .ip1(\pipeline/regfile/data[4][25] ), .ip2(n18344), .s(
        n19383), .op(n9775) );
  nand2_1 U20573 ( .ip1(\pipeline/PC_IF [26]), .ip2(n21996), .op(n18345) );
  nand2_1 U20574 ( .ip1(n18346), .ip2(n18345), .op(n8438) );
  nand2_1 U20575 ( .ip1(\pipeline/PC_IF [26]), .ip2(n21988), .op(n18348) );
  nand2_1 U20576 ( .ip1(\pipeline/PC_DX [26]), .ip2(n21999), .op(n18347) );
  nand2_1 U20577 ( .ip1(n18348), .ip2(n18347), .op(n8437) );
  nand2_1 U20578 ( .ip1(n18350), .ip2(n18349), .op(n18359) );
  inv_1 U20579 ( .ip(n18351), .op(n18725) );
  nor2_1 U20580 ( .ip1(n18354), .ip2(n18725), .op(n18352) );
  nor2_1 U20581 ( .ip1(n18353), .ip2(n18352), .op(n18357) );
  inv_1 U20582 ( .ip(n18354), .op(n18722) );
  nand2_1 U20583 ( .ip1(n18723), .ip2(n18722), .op(n18355) );
  or2_1 U20584 ( .ip1(n18355), .ip2(n19177), .op(n18356) );
  nand2_1 U20585 ( .ip1(n18357), .ip2(n18356), .op(n18358) );
  xnor2_1 U20586 ( .ip1(n18359), .ip2(n18358), .op(n18360) );
  nand2_1 U20587 ( .ip1(n18360), .ip2(n21577), .op(n18385) );
  nand4_1 U20588 ( .ip1(n18364), .ip2(n18363), .ip3(n18362), .ip4(n18361), 
        .op(n18937) );
  nand2_1 U20589 ( .ip1(n18937), .ip2(n19427), .op(n18366) );
  nand2_1 U20590 ( .ip1(n18935), .ip2(n21540), .op(n18365) );
  nand2_1 U20591 ( .ip1(n18366), .ip2(n18365), .op(n18381) );
  nand2_1 U20592 ( .ip1(n18934), .ip2(n18367), .op(n18377) );
  nor3_1 U20593 ( .ip1(n18368), .ip2(n21551), .ip3(n11941), .op(n18372) );
  nor2_1 U20594 ( .ip1(n18369), .ip2(n16914), .op(n18370) );
  nor2_1 U20595 ( .ip1(n20907), .ip2(n18370), .op(n18371) );
  not_ab_or_c_or_d U20596 ( .ip1(n20911), .ip2(n18373), .ip3(n18372), .ip4(
        n18371), .op(n18376) );
  nand2_1 U20597 ( .ip1(n18944), .ip2(n18374), .op(n18375) );
  nor2_1 U20598 ( .ip1(n20883), .ip2(n18378), .op(n18379) );
  not_ab_or_c_or_d U20599 ( .ip1(n20900), .ip2(n18381), .ip3(n18380), .ip4(
        n18379), .op(n18384) );
  nand2_1 U20600 ( .ip1(n18382), .ip2(n13166), .op(n18383) );
  nand3_1 U20601 ( .ip1(n18385), .ip2(n18384), .ip3(n18383), .op(
        dmem_haddr[25]) );
  mux2_1 U20602 ( .ip1(dmem_haddr[25]), .ip2(\pipeline/alu_out_WB [25]), .s(
        n19505), .op(n8707) );
  nand2_1 U20603 ( .ip1(\pipeline/ctrl/prev_ex_code_WB [0]), .ip2(n19505), 
        .op(n18393) );
  nor2_1 U20604 ( .ip1(\pipeline/ctrl/had_ex_DX ), .ip2(n19505), .op(n21099)
         );
  nand3_1 U20605 ( .ip1(\pipeline/prv [0]), .ip2(n21095), .ip3(n21097), .op(
        n18390) );
  inv_1 U20606 ( .ip(n18386), .op(n18387) );
  nand2_1 U20607 ( .ip1(n18388), .ip2(n18387), .op(n18389) );
  nand2_1 U20608 ( .ip1(n18390), .ip2(n18389), .op(n18391) );
  nand2_1 U20609 ( .ip1(n21099), .ip2(n18391), .op(n18392) );
  nand2_1 U20610 ( .ip1(n18393), .ip2(n18392), .op(n8738) );
  nand2_1 U20611 ( .ip1(\pipeline/ctrl/prev_ex_code_WB [3]), .ip2(n19505), 
        .op(n18395) );
  nand3_1 U20612 ( .ip1(n21095), .ip2(n21097), .ip3(n21099), .op(n18394) );
  nand2_1 U20613 ( .ip1(n18395), .ip2(n18394), .op(n8739) );
  inv_1 U20614 ( .ip(n21110), .op(n20844) );
  nand2_1 U20615 ( .ip1(n20844), .ip2(n19677), .op(n18399) );
  nand2_1 U20616 ( .ip1(\pipeline/csr/instret_full [39]), .ip2(n21117), .op(
        n18398) );
  inv_1 U20617 ( .ip(n21111), .op(n20334) );
  or2_1 U20618 ( .ip1(\pipeline/csr/instret_full [39]), .ip2(n20338), .op(
        n18396) );
  nand3_1 U20619 ( .ip1(n18400), .ip2(n20334), .ip3(n18396), .op(n18397) );
  nand3_1 U20620 ( .ip1(n18399), .ip2(n18398), .ip3(n18397), .op(n10099) );
  nor2_1 U20621 ( .ip1(n19700), .ip2(n21110), .op(n18403) );
  not_ab_or_c_or_d U20622 ( .ip1(n18401), .ip2(n18400), .ip3(n21111), .ip4(
        n18471), .op(n18402) );
  ab_or_c_or_d U20623 ( .ip1(n21117), .ip2(\pipeline/csr/instret_full [40]), 
        .ip3(n18403), .ip4(n18402), .op(n10098) );
  nand2_1 U20624 ( .ip1(n21032), .ip2(n18470), .op(n18405) );
  nand2_1 U20625 ( .ip1(\pipeline/csr/mtvec [9]), .ip2(n20705), .op(n18404) );
  nand2_1 U20626 ( .ip1(n18405), .ip2(n18404), .op(n9983) );
  nand2_1 U20627 ( .ip1(\pipeline/csr/from_host [9]), .ip2(n22372), .op(n18407) );
  nand2_1 U20628 ( .ip1(n22373), .ip2(n18470), .op(n18406) );
  nand2_1 U20629 ( .ip1(n18407), .ip2(n18406), .op(n9951) );
  nand2_1 U20630 ( .ip1(n22378), .ip2(n18470), .op(n18409) );
  nand2_1 U20631 ( .ip1(\pipeline/csr/to_host [9]), .ip2(n22376), .op(n18408)
         );
  nand2_1 U20632 ( .ip1(n18409), .ip2(n18408), .op(n8763) );
  inv_1 U20633 ( .ip(\pipeline/csr/instret_full [9]), .op(n18411) );
  nor2_1 U20634 ( .ip1(n18411), .ip2(n20990), .op(n18414) );
  mux2_1 U20635 ( .ip1(n18411), .ip2(\pipeline/csr/instret_full [9]), .s(
        n18410), .op(n18412) );
  nor2_1 U20636 ( .ip1(n21005), .ip2(n18412), .op(n18413) );
  ab_or_c_or_d U20637 ( .ip1(n21019), .ip2(n18470), .ip3(n18414), .ip4(n18413), 
        .op(n10129) );
  inv_1 U20638 ( .ip(n18470), .op(n18466) );
  nor2_1 U20639 ( .ip1(n18466), .ip2(n21168), .op(n18417) );
  xor2_1 U20640 ( .ip1(\pipeline/PC_WB [9]), .ip2(n19771), .op(n18415) );
  nor2_1 U20641 ( .ip1(n21171), .ip2(n18415), .op(n18416) );
  ab_or_c_or_d U20642 ( .ip1(n21174), .ip2(\pipeline/epc [9]), .ip3(n18417), 
        .ip4(n18416), .op(n8862) );
  nand2_1 U20643 ( .ip1(n21238), .ip2(dmem_rdata[9]), .op(n18418) );
  or2_1 U20644 ( .ip1(n18418), .ip2(n22071), .op(n18421) );
  nand2_1 U20645 ( .ip1(n19386), .ip2(dmem_rdata[17]), .op(n18419) );
  or2_1 U20646 ( .ip1(n18419), .ip2(n22071), .op(n18420) );
  nand2_1 U20647 ( .ip1(n18421), .ip2(n18420), .op(n18422) );
  not_ab_or_c_or_d U20648 ( .ip1(n18423), .ip2(n21583), .ip3(n18422), .ip4(
        n19390), .op(n18426) );
  inv_1 U20649 ( .ip(n21240), .op(n18424) );
  nor2_1 U20650 ( .ip1(n22071), .ip2(n18424), .op(n19410) );
  nand2_1 U20651 ( .ip1(dmem_rdata[25]), .ip2(n19410), .op(n18425) );
  nand2_1 U20652 ( .ip1(n18426), .ip2(n18425), .op(n18427) );
  mux2_1 U20653 ( .ip1(\pipeline/regfile/data[29][9] ), .ip2(n18427), .s(
        n21619), .op(n8991) );
  mux2_1 U20654 ( .ip1(\pipeline/regfile/data[14][9] ), .ip2(n18427), .s(
        n21604), .op(n9471) );
  mux2_1 U20655 ( .ip1(\pipeline/regfile/data[22][9] ), .ip2(n18427), .s(
        n21589), .op(n9215) );
  mux2_1 U20656 ( .ip1(\pipeline/regfile/data[5][9] ), .ip2(n18427), .s(n21598), .op(n9759) );
  mux2_1 U20657 ( .ip1(\pipeline/regfile/data[27][9] ), .ip2(n18427), .s(
        n21612), .op(n9055) );
  mux2_1 U20658 ( .ip1(\pipeline/regfile/data[26][9] ), .ip2(n18427), .s(
        n21607), .op(n9087) );
  mux2_1 U20659 ( .ip1(\pipeline/regfile/data[28][9] ), .ip2(n18427), .s(
        n21590), .op(n9023) );
  mux2_1 U20660 ( .ip1(\pipeline/regfile/data[31][9] ), .ip2(n18427), .s(
        n21606), .op(n8927) );
  mux2_1 U20661 ( .ip1(\pipeline/regfile/data[19][9] ), .ip2(n18427), .s(
        n21592), .op(n9311) );
  mux2_1 U20662 ( .ip1(\pipeline/regfile/data[6][9] ), .ip2(n18427), .s(n21597), .op(n9727) );
  mux2_1 U20663 ( .ip1(\pipeline/regfile/data[30][9] ), .ip2(n18427), .s(
        n21594), .op(n8959) );
  mux2_1 U20664 ( .ip1(\pipeline/regfile/data[18][9] ), .ip2(n18427), .s(
        n21595), .op(n9343) );
  mux2_1 U20665 ( .ip1(\pipeline/regfile/data[11][9] ), .ip2(n18427), .s(
        n21593), .op(n9567) );
  mux2_1 U20666 ( .ip1(\pipeline/regfile/data[25][9] ), .ip2(n18427), .s(
        n21602), .op(n9119) );
  mux2_1 U20667 ( .ip1(\pipeline/regfile/data[13][9] ), .ip2(n18427), .s(
        n21600), .op(n9503) );
  mux2_1 U20668 ( .ip1(\pipeline/regfile/data[17][9] ), .ip2(n18427), .s(
        n21616), .op(n9375) );
  mux2_1 U20669 ( .ip1(\pipeline/regfile/data[23][9] ), .ip2(n18427), .s(
        n21596), .op(n9183) );
  mux2_1 U20670 ( .ip1(\pipeline/regfile/data[12][9] ), .ip2(n18427), .s(
        n21591), .op(n9535) );
  mux2_1 U20671 ( .ip1(\pipeline/regfile/data[7][9] ), .ip2(n18427), .s(n21614), .op(n9695) );
  mux2_1 U20672 ( .ip1(\pipeline/regfile/data[8][9] ), .ip2(n18427), .s(n21617), .op(n9663) );
  mux2_1 U20673 ( .ip1(\pipeline/regfile/data[15][9] ), .ip2(n18427), .s(
        n21613), .op(n9439) );
  mux2_1 U20674 ( .ip1(\pipeline/regfile/data[10][9] ), .ip2(n18427), .s(
        n21618), .op(n9599) );
  mux2_1 U20675 ( .ip1(\pipeline/regfile/data[21][9] ), .ip2(n18427), .s(
        n21615), .op(n9247) );
  mux2_1 U20676 ( .ip1(\pipeline/regfile/data[24][9] ), .ip2(n18427), .s(
        n21603), .op(n9151) );
  mux2_1 U20677 ( .ip1(\pipeline/regfile/data[20][9] ), .ip2(n18427), .s(
        n21601), .op(n9279) );
  mux2_1 U20678 ( .ip1(\pipeline/regfile/data[9][9] ), .ip2(n18427), .s(n21609), .op(n9631) );
  mux2_1 U20679 ( .ip1(\pipeline/regfile/data[16][9] ), .ip2(n18427), .s(
        n21608), .op(n9407) );
  mux2_1 U20680 ( .ip1(\pipeline/regfile/data[3][9] ), .ip2(n18427), .s(n21599), .op(n9823) );
  mux2_1 U20681 ( .ip1(\pipeline/regfile/data[1][9] ), .ip2(n18427), .s(n21611), .op(n9887) );
  mux2_1 U20682 ( .ip1(\pipeline/regfile/data[2][9] ), .ip2(n18427), .s(n21610), .op(n9855) );
  mux2_1 U20683 ( .ip1(\pipeline/regfile/data[4][9] ), .ip2(n18427), .s(n21605), .op(n9791) );
  mux2_1 U20684 ( .ip1(dmem_haddr[9]), .ip2(\pipeline/alu_out_WB [9]), .s(
        n21582), .op(n8723) );
  inv_1 U20685 ( .ip(n18428), .op(n18429) );
  nor2_1 U20686 ( .ip1(\pipeline/csr/time_full [9]), .ip2(n18429), .op(n18431)
         );
  nor3_1 U20687 ( .ip1(n21177), .ip2(n19784), .ip3(n18431), .op(n18430) );
  not_ab_or_c_or_d U20688 ( .ip1(n21179), .ip2(n18470), .ip3(n21217), .ip4(
        n18430), .op(n18434) );
  buf_1 U20689 ( .ip(n21198), .op(n22254) );
  nor2_1 U20690 ( .ip1(n18431), .ip2(n19784), .op(n18432) );
  nor2_1 U20691 ( .ip1(n22254), .ip2(n18432), .op(n18433) );
  nor2_1 U20692 ( .ip1(n18434), .ip2(n18433), .op(\pipeline/csr/N1946 ) );
  inv_1 U20693 ( .ip(n18435), .op(n20748) );
  nor2_1 U20694 ( .ip1(n20748), .ip2(n21210), .op(n22282) );
  inv_1 U20695 ( .ip(n22282), .op(n22267) );
  nor2_1 U20696 ( .ip1(n18466), .ip2(n22267), .op(n18438) );
  not_ab_or_c_or_d U20697 ( .ip1(n19697), .ip2(n18436), .ip3(n19780), .ip4(
        n22276), .op(n18437) );
  or2_1 U20698 ( .ip1(n18438), .ip2(n18437), .op(\pipeline/csr/N1978 ) );
  or3_1 U20699 ( .ip1(\pipeline/inst_DX [26]), .ip2(n21089), .ip3(n18439), 
        .op(n18446) );
  inv_1 U20700 ( .ip(n18446), .op(n21195) );
  nand2_1 U20701 ( .ip1(n21198), .ip2(n21195), .op(n21131) );
  inv_1 U20702 ( .ip(n21131), .op(n22008) );
  nand2_1 U20703 ( .ip1(n22008), .ip2(n18470), .op(n18443) );
  inv_1 U20704 ( .ip(\pipeline/csr/mtime_full [4]), .op(n19622) );
  inv_1 U20705 ( .ip(\pipeline/csr/mtime_full [2]), .op(n19623) );
  inv_1 U20706 ( .ip(\pipeline/csr/mtime_full [1]), .op(n19635) );
  inv_1 U20707 ( .ip(\pipeline/csr/mtime_full [0]), .op(n20980) );
  nor3_1 U20708 ( .ip1(n19623), .ip2(n19635), .ip3(n20980), .op(n21192) );
  nand2_1 U20709 ( .ip1(\pipeline/csr/mtime_full [3]), .ip2(n21192), .op(
        n20820) );
  nor2_1 U20710 ( .ip1(n19622), .ip2(n20820), .op(n21063) );
  nand2_1 U20711 ( .ip1(\pipeline/csr/mtime_full [5]), .ip2(n21063), .op(
        n20350) );
  nor2_1 U20712 ( .ip1(n19659), .ip2(n20350), .op(n20353) );
  nand2_1 U20713 ( .ip1(\pipeline/csr/mtime_full [7]), .ip2(n20353), .op(
        n19708) );
  nor2_1 U20714 ( .ip1(n19637), .ip2(n19708), .op(n19711) );
  xor2_1 U20715 ( .ip1(\pipeline/csr/mtime_full [9]), .ip2(n19711), .op(n18441) );
  nand2_1 U20716 ( .ip1(n20966), .ip2(n18439), .op(n18447) );
  or2_1 U20717 ( .ip1(htif_reset), .ip2(n18440), .op(n19804) );
  nand2_1 U20718 ( .ip1(n18447), .ip2(n19804), .op(n18532) );
  nor2_1 U20719 ( .ip1(n21120), .ip2(n18532), .op(n21134) );
  inv_1 U20720 ( .ip(n21134), .op(n22009) );
  nand2_1 U20721 ( .ip1(n18441), .ip2(n22009), .op(n18442) );
  nand2_1 U20722 ( .ip1(n18443), .ip2(n18442), .op(\pipeline/csr/N2090 ) );
  nand2_1 U20723 ( .ip1(\pipeline/csr/mscratch [9]), .ip2(n22013), .op(n18445)
         );
  nand2_1 U20724 ( .ip1(n22014), .ip2(n18470), .op(n18444) );
  nand2_1 U20725 ( .ip1(n18445), .ip2(n18444), .op(n9919) );
  nand2_1 U20726 ( .ip1(n18447), .ip2(n18446), .op(n18448) );
  or2_1 U20727 ( .ip1(n18448), .ip2(n21120), .op(n18449) );
  inv_1 U20728 ( .ip(\pipeline/csr/mtime_full [36]), .op(n22142) );
  inv_1 U20729 ( .ip(\pipeline/csr/mtime_full [34]), .op(n22137) );
  inv_1 U20730 ( .ip(\pipeline/csr/mtime_full [32]), .op(n22125) );
  inv_1 U20731 ( .ip(\pipeline/csr/mtime_full [30]), .op(n19638) );
  inv_1 U20732 ( .ip(\pipeline/csr/mtime_full [28]), .op(n19620) );
  inv_1 U20733 ( .ip(\pipeline/csr/mtime_full [26]), .op(n19660) );
  inv_1 U20734 ( .ip(\pipeline/csr/mtime_full [24]), .op(n19621) );
  inv_1 U20735 ( .ip(\pipeline/csr/mtime_full [22]), .op(n19604) );
  inv_1 U20736 ( .ip(\pipeline/csr/mtime_full [18]), .op(n19610) );
  inv_1 U20737 ( .ip(\pipeline/csr/mtime_full [16]), .op(n19629) );
  inv_1 U20738 ( .ip(\pipeline/csr/mtime_full [14]), .op(n19650) );
  inv_1 U20739 ( .ip(\pipeline/csr/mtime_full [12]), .op(n19630) );
  inv_1 U20740 ( .ip(\pipeline/csr/mtime_full [10]), .op(n19636) );
  nand2_1 U20741 ( .ip1(\pipeline/csr/mtime_full [9]), .ip2(n19711), .op(
        n19791) );
  nor2_1 U20742 ( .ip1(n19636), .ip2(n19791), .op(n20168) );
  nand2_1 U20743 ( .ip1(\pipeline/csr/mtime_full [11]), .ip2(n20168), .op(
        n20758) );
  nor2_1 U20744 ( .ip1(n19630), .ip2(n20758), .op(n20761) );
  nand2_1 U20745 ( .ip1(\pipeline/csr/mtime_full [13]), .ip2(n20761), .op(
        n19857) );
  nor2_1 U20746 ( .ip1(n19650), .ip2(n19857), .op(n19860) );
  nand2_1 U20747 ( .ip1(\pipeline/csr/mtime_full [15]), .ip2(n19860), .op(
        n19914) );
  nor2_1 U20748 ( .ip1(n19629), .ip2(n19914), .op(n19966) );
  nand2_1 U20749 ( .ip1(\pipeline/csr/mtime_full [17]), .ip2(n19966), .op(
        n18530) );
  nor2_1 U20750 ( .ip1(n19610), .ip2(n18530), .op(n18595) );
  nand2_1 U20751 ( .ip1(\pipeline/csr/mtime_full [19]), .ip2(n18595), .op(
        n19518) );
  nor2_1 U20752 ( .ip1(n19658), .ip2(n19518), .op(n19521) );
  nand2_1 U20753 ( .ip1(\pipeline/csr/mtime_full [21]), .ip2(n19521), .op(
        n20070) );
  nor2_1 U20754 ( .ip1(n19604), .ip2(n20070), .op(n20123) );
  nand2_1 U20755 ( .ip1(\pipeline/csr/mtime_full [23]), .ip2(n20123), .op(
        n18761) );
  nor2_1 U20756 ( .ip1(n19621), .ip2(n18761), .op(n18807) );
  nand2_1 U20757 ( .ip1(\pipeline/csr/mtime_full [25]), .ip2(n18807), .op(
        n19102) );
  nor2_1 U20758 ( .ip1(n19660), .ip2(n19102), .op(n19155) );
  nand2_1 U20759 ( .ip1(\pipeline/csr/mtime_full [27]), .ip2(n19155), .op(
        n19262) );
  nor2_1 U20760 ( .ip1(n19620), .ip2(n19262), .op(n19265) );
  nand2_1 U20761 ( .ip1(\pipeline/csr/mtime_full [29]), .ip2(n19265), .op(
        n18985) );
  nor2_1 U20762 ( .ip1(n19638), .ip2(n18985), .op(n20935) );
  nand2_1 U20763 ( .ip1(\pipeline/csr/mtime_full [31]), .ip2(n20935), .op(
        n22124) );
  nor2_1 U20764 ( .ip1(n22125), .ip2(n22124), .op(n22130) );
  nand2_1 U20765 ( .ip1(\pipeline/csr/mtime_full [33]), .ip2(n22130), .op(
        n22136) );
  nor2_1 U20766 ( .ip1(n22137), .ip2(n22136), .op(n22135) );
  nand2_1 U20767 ( .ip1(\pipeline/csr/mtime_full [35]), .ip2(n22135), .op(
        n22141) );
  nor2_1 U20768 ( .ip1(n22142), .ip2(n22141), .op(n22146) );
  nand2_1 U20769 ( .ip1(\pipeline/csr/mtime_full [37]), .ip2(n22146), .op(
        n22152) );
  nor2_1 U20770 ( .ip1(n22153), .ip2(n22152), .op(n22151) );
  nand2_1 U20771 ( .ip1(\pipeline/csr/mtime_full [39]), .ip2(n22151), .op(
        n19723) );
  nor2_1 U20772 ( .ip1(n18450), .ip2(n19723), .op(n19722) );
  xor2_1 U20773 ( .ip1(\pipeline/csr/mtime_full [41]), .ip2(n19722), .op(
        n18451) );
  nand2_1 U20774 ( .ip1(n18449), .ip2(n18451), .op(n18454) );
  inv_1 U20775 ( .ip(n19804), .op(n21208) );
  nand2_1 U20776 ( .ip1(n21208), .ip2(n18470), .op(n18452) );
  or2_1 U20777 ( .ip1(n21210), .ip2(n18452), .op(n18453) );
  nand2_1 U20778 ( .ip1(n18454), .ip2(n18453), .op(\pipeline/csr/N2122 ) );
  or2_1 U20779 ( .ip1(n21089), .ip2(n18456), .op(n18605) );
  inv_1 U20780 ( .ip(n19731), .op(n18455) );
  nor2_1 U20781 ( .ip1(\pipeline/csr/cycle_full [9]), .ip2(n18455), .op(n18458) );
  nand2_1 U20782 ( .ip1(n20966), .ip2(n18456), .op(n21215) );
  nor3_1 U20783 ( .ip1(n19811), .ip2(n18458), .ip3(n21215), .op(n18457) );
  not_ab_or_c_or_d U20784 ( .ip1(n21076), .ip2(n18470), .ip3(n21120), .ip4(
        n18457), .op(n18461) );
  nor2_1 U20785 ( .ip1(n18458), .ip2(n19811), .op(n18459) );
  nor2_1 U20786 ( .ip1(n22254), .ip2(n18459), .op(n18460) );
  nor2_1 U20787 ( .ip1(n18461), .ip2(n18460), .op(\pipeline/csr/N1882 ) );
  nand2_1 U20788 ( .ip1(\pipeline/csr/mtimecmp [9]), .ip2(n22363), .op(n18463)
         );
  nand2_1 U20789 ( .ip1(n22365), .ip2(n18470), .op(n18462) );
  nand2_1 U20790 ( .ip1(n18463), .ip2(n18462), .op(n10013) );
  nand2_1 U20791 ( .ip1(\pipeline/csr/mie [9]), .ip2(n22356), .op(n18465) );
  nand2_1 U20792 ( .ip1(n22357), .ip2(n18470), .op(n18464) );
  nand2_1 U20793 ( .ip1(n18465), .ip2(n18464), .op(n10051) );
  nor2_1 U20794 ( .ip1(n18466), .ip2(n22305), .op(n18469) );
  not_ab_or_c_or_d U20795 ( .ip1(n19742), .ip2(n18467), .ip3(n19829), .ip4(
        n22308), .op(n18468) );
  or2_1 U20796 ( .ip1(n18469), .ip2(n18468), .op(\pipeline/csr/N1914 ) );
  nand2_1 U20797 ( .ip1(n20844), .ip2(n18470), .op(n18475) );
  nand2_1 U20798 ( .ip1(\pipeline/csr/instret_full [41]), .ip2(n21117), .op(
        n18474) );
  or2_1 U20799 ( .ip1(\pipeline/csr/instret_full [41]), .ip2(n18471), .op(
        n18472) );
  nand3_1 U20800 ( .ip1(n18477), .ip2(n20334), .ip3(n18472), .op(n18473) );
  nand3_1 U20801 ( .ip1(n18475), .ip2(n18474), .ip3(n18473), .op(n10097) );
  nor2_1 U20802 ( .ip1(n19805), .ip2(n21110), .op(n18480) );
  not_ab_or_c_or_d U20803 ( .ip1(n18478), .ip2(n18477), .ip3(n21111), .ip4(
        n18476), .op(n18479) );
  ab_or_c_or_d U20804 ( .ip1(n21117), .ip2(\pipeline/csr/instret_full [42]), 
        .ip3(n18480), .ip4(n18479), .op(n10096) );
  nand2_1 U20805 ( .ip1(n20788), .ip2(n20844), .op(n18486) );
  and2_1 U20806 ( .ip1(n21117), .ip2(\pipeline/csr/instret_full [44]), .op(
        n18484) );
  inv_1 U20807 ( .ip(\pipeline/csr/instret_full [44]), .op(n18482) );
  nor2_1 U20808 ( .ip1(n18482), .ip2(n18481), .op(n18487) );
  not_ab_or_c_or_d U20809 ( .ip1(n18482), .ip2(n18481), .ip3(n18487), .ip4(
        n21111), .op(n18483) );
  nor2_1 U20810 ( .ip1(n18484), .ip2(n18483), .op(n18485) );
  nand2_1 U20811 ( .ip1(n18486), .ip2(n18485), .op(n10094) );
  nand2_1 U20812 ( .ip1(n20844), .ip2(n22166), .op(n18491) );
  nand2_1 U20813 ( .ip1(\pipeline/csr/instret_full [45]), .ip2(n21117), .op(
        n18490) );
  nand2_1 U20814 ( .ip1(\pipeline/csr/instret_full [45]), .ip2(n18487), .op(
        n18492) );
  or2_1 U20815 ( .ip1(\pipeline/csr/instret_full [45]), .ip2(n18487), .op(
        n18488) );
  nand3_1 U20816 ( .ip1(n18492), .ip2(n20334), .ip3(n18488), .op(n18489) );
  nand3_1 U20817 ( .ip1(n18491), .ip2(n18490), .ip3(n18489), .op(n10093) );
  inv_1 U20818 ( .ip(\pipeline/csr/instret_full [46]), .op(n18493) );
  nor2_1 U20819 ( .ip1(n18493), .ip2(n18492), .op(n18496) );
  not_ab_or_c_or_d U20820 ( .ip1(n18493), .ip2(n18492), .ip3(n21111), .ip4(
        n18496), .op(n18495) );
  nor2_1 U20821 ( .ip1(n18493), .ip2(n19134), .op(n18494) );
  ab_or_c_or_d U20822 ( .ip1(n20844), .ip2(n22171), .ip3(n18495), .ip4(n18494), 
        .op(n10092) );
  nand2_1 U20823 ( .ip1(n20844), .ip2(n22177), .op(n18500) );
  nand2_1 U20824 ( .ip1(\pipeline/csr/instret_full [47]), .ip2(n21117), .op(
        n18499) );
  nand2_1 U20825 ( .ip1(\pipeline/csr/instret_full [47]), .ip2(n18496), .op(
        n18501) );
  or2_1 U20826 ( .ip1(\pipeline/csr/instret_full [47]), .ip2(n18496), .op(
        n18497) );
  nand3_1 U20827 ( .ip1(n18501), .ip2(n20334), .ip3(n18497), .op(n18498) );
  nand3_1 U20828 ( .ip1(n18500), .ip2(n18499), .ip3(n18498), .op(n10091) );
  inv_1 U20829 ( .ip(\pipeline/csr/instret_full [48]), .op(n18502) );
  nor2_1 U20830 ( .ip1(n18502), .ip2(n18501), .op(n18505) );
  not_ab_or_c_or_d U20831 ( .ip1(n18502), .ip2(n18501), .ip3(n21111), .ip4(
        n18505), .op(n18504) );
  inv_1 U20832 ( .ip(n21117), .op(n19134) );
  nor2_1 U20833 ( .ip1(n18502), .ip2(n19134), .op(n18503) );
  ab_or_c_or_d U20834 ( .ip1(n20844), .ip2(n19951), .ip3(n18504), .ip4(n18503), 
        .op(n10090) );
  nand2_1 U20835 ( .ip1(n20844), .ip2(n22183), .op(n18509) );
  nand2_1 U20836 ( .ip1(\pipeline/csr/instret_full [49]), .ip2(n21117), .op(
        n18508) );
  nand2_1 U20837 ( .ip1(\pipeline/csr/instret_full [49]), .ip2(n18505), .op(
        n18573) );
  or2_1 U20838 ( .ip1(\pipeline/csr/instret_full [49]), .ip2(n18505), .op(
        n18506) );
  nand3_1 U20839 ( .ip1(n18573), .ip2(n20334), .ip3(n18506), .op(n18507) );
  nand3_1 U20840 ( .ip1(n18509), .ip2(n18508), .ip3(n18507), .op(n10089) );
  nor2_1 U20841 ( .ip1(n18572), .ip2(n21168), .op(n18512) );
  xor2_1 U20842 ( .ip1(\pipeline/PC_WB [18]), .ip2(n20028), .op(n18510) );
  nor2_1 U20843 ( .ip1(n21171), .ip2(n18510), .op(n18511) );
  ab_or_c_or_d U20844 ( .ip1(n21174), .ip2(\pipeline/epc [18]), .ip3(n18512), 
        .ip4(n18511), .op(n8853) );
  nand2_1 U20845 ( .ip1(n21032), .ip2(n18563), .op(n18514) );
  nand2_1 U20846 ( .ip1(\pipeline/csr/mtvec [18]), .ip2(n20705), .op(n18513)
         );
  nand2_1 U20847 ( .ip1(n18514), .ip2(n18513), .op(n9974) );
  nand2_1 U20848 ( .ip1(n21585), .ip2(dmem_rdata[18]), .op(n18519) );
  nand2_1 U20849 ( .ip1(n18515), .ip2(n21583), .op(n18518) );
  nor2_1 U20850 ( .ip1(n18516), .ip2(n19302), .op(n19324) );
  nand2_1 U20851 ( .ip1(dmem_rdata[26]), .ip2(n19324), .op(n18517) );
  nand4_1 U20852 ( .ip1(n21588), .ip2(n18519), .ip3(n18518), .ip4(n18517), 
        .op(n18520) );
  mux2_1 U20853 ( .ip1(\pipeline/regfile/data[29][18] ), .ip2(n18520), .s(
        n19353), .op(n8982) );
  mux2_1 U20854 ( .ip1(\pipeline/regfile/data[14][18] ), .ip2(n18520), .s(
        n19354), .op(n9462) );
  mux2_1 U20855 ( .ip1(\pipeline/regfile/data[22][18] ), .ip2(n18520), .s(
        n19355), .op(n9206) );
  mux2_1 U20856 ( .ip1(\pipeline/regfile/data[5][18] ), .ip2(n18520), .s(
        n19356), .op(n9750) );
  mux2_1 U20857 ( .ip1(\pipeline/regfile/data[27][18] ), .ip2(n18520), .s(
        n19357), .op(n9046) );
  mux2_1 U20858 ( .ip1(\pipeline/regfile/data[26][18] ), .ip2(n18520), .s(
        n19358), .op(n9078) );
  mux2_1 U20859 ( .ip1(\pipeline/regfile/data[28][18] ), .ip2(n18520), .s(
        n19359), .op(n9014) );
  mux2_1 U20860 ( .ip1(\pipeline/regfile/data[31][18] ), .ip2(n18520), .s(
        n19360), .op(n8918) );
  mux2_1 U20861 ( .ip1(\pipeline/regfile/data[19][18] ), .ip2(n18520), .s(
        n19361), .op(n9302) );
  mux2_1 U20862 ( .ip1(\pipeline/regfile/data[6][18] ), .ip2(n18520), .s(
        n19362), .op(n9718) );
  mux2_1 U20863 ( .ip1(\pipeline/regfile/data[30][18] ), .ip2(n18520), .s(
        n19363), .op(n8950) );
  mux2_1 U20864 ( .ip1(\pipeline/regfile/data[18][18] ), .ip2(n18520), .s(
        n19364), .op(n9334) );
  mux2_1 U20865 ( .ip1(\pipeline/regfile/data[11][18] ), .ip2(n18520), .s(
        n19365), .op(n9558) );
  mux2_1 U20866 ( .ip1(\pipeline/regfile/data[25][18] ), .ip2(n18520), .s(
        n19366), .op(n9110) );
  mux2_1 U20867 ( .ip1(\pipeline/regfile/data[13][18] ), .ip2(n18520), .s(
        n19367), .op(n9494) );
  mux2_1 U20868 ( .ip1(\pipeline/regfile/data[17][18] ), .ip2(n18520), .s(
        n19368), .op(n9366) );
  mux2_1 U20869 ( .ip1(\pipeline/regfile/data[23][18] ), .ip2(n18520), .s(
        n19369), .op(n9174) );
  mux2_1 U20870 ( .ip1(\pipeline/regfile/data[12][18] ), .ip2(n18520), .s(
        n19370), .op(n9526) );
  mux2_1 U20871 ( .ip1(\pipeline/regfile/data[7][18] ), .ip2(n18520), .s(
        n19371), .op(n9686) );
  mux2_1 U20872 ( .ip1(\pipeline/regfile/data[8][18] ), .ip2(n18520), .s(
        n19372), .op(n9654) );
  mux2_1 U20873 ( .ip1(\pipeline/regfile/data[15][18] ), .ip2(n18520), .s(
        n19373), .op(n9430) );
  mux2_1 U20874 ( .ip1(\pipeline/regfile/data[10][18] ), .ip2(n18520), .s(
        n19374), .op(n9590) );
  mux2_1 U20875 ( .ip1(\pipeline/regfile/data[21][18] ), .ip2(n18520), .s(
        n19375), .op(n9238) );
  mux2_1 U20876 ( .ip1(\pipeline/regfile/data[24][18] ), .ip2(n18520), .s(
        n19376), .op(n9142) );
  mux2_1 U20877 ( .ip1(\pipeline/regfile/data[20][18] ), .ip2(n18520), .s(
        n19377), .op(n9270) );
  mux2_1 U20878 ( .ip1(\pipeline/regfile/data[9][18] ), .ip2(n18520), .s(
        n19378), .op(n9622) );
  mux2_1 U20879 ( .ip1(\pipeline/regfile/data[16][18] ), .ip2(n18520), .s(
        n19379), .op(n9398) );
  mux2_1 U20880 ( .ip1(\pipeline/regfile/data[3][18] ), .ip2(n18520), .s(
        n19380), .op(n9814) );
  mux2_1 U20881 ( .ip1(\pipeline/regfile/data[1][18] ), .ip2(n18520), .s(
        n19381), .op(n9878) );
  mux2_1 U20882 ( .ip1(\pipeline/regfile/data[2][18] ), .ip2(n18520), .s(
        n19382), .op(n9846) );
  mux2_1 U20883 ( .ip1(\pipeline/regfile/data[4][18] ), .ip2(n18520), .s(
        n19383), .op(n9782) );
  mux2_1 U20884 ( .ip1(dmem_haddr[18]), .ip2(\pipeline/alu_out_WB [18]), .s(
        n21582), .op(n8714) );
  or2_1 U20885 ( .ip1(\pipeline/csr/time_full [50]), .ip2(n19972), .op(n18521)
         );
  nand2_1 U20886 ( .ip1(n18585), .ip2(n18521), .op(n18522) );
  or2_1 U20887 ( .ip1(n22276), .ip2(n18522), .op(n18524) );
  nand2_1 U20888 ( .ip1(n22282), .ip2(n18563), .op(n18523) );
  nand2_1 U20889 ( .ip1(n18524), .ip2(n18523), .op(\pipeline/csr/N1987 ) );
  nor2_1 U20890 ( .ip1(n22252), .ip2(n21120), .op(n22002) );
  or2_1 U20891 ( .ip1(\pipeline/csr/time_full [18]), .ip2(n19980), .op(n18525)
         );
  nand2_1 U20892 ( .ip1(n18588), .ip2(n18525), .op(n18526) );
  or2_1 U20893 ( .ip1(n22002), .ip2(n18526), .op(n18529) );
  inv_1 U20894 ( .ip(n21179), .op(n18527) );
  nor2_1 U20895 ( .ip1(n18527), .ip2(n21210), .op(n22005) );
  nand2_1 U20896 ( .ip1(n22005), .ip2(n18563), .op(n18528) );
  nand2_1 U20897 ( .ip1(n18529), .ip2(n18528), .op(\pipeline/csr/N1955 ) );
  inv_1 U20898 ( .ip(n18530), .op(n18531) );
  nor2_1 U20899 ( .ip1(\pipeline/csr/mtime_full [18]), .ip2(n18531), .op(
        n18534) );
  inv_1 U20900 ( .ip(n18532), .op(n21193) );
  nor3_1 U20901 ( .ip1(n18534), .ip2(n21193), .ip3(n18595), .op(n18533) );
  not_ab_or_c_or_d U20902 ( .ip1(n21195), .ip2(n18563), .ip3(n21120), .ip4(
        n18533), .op(n18537) );
  nor2_1 U20903 ( .ip1(n18534), .ip2(n18595), .op(n18535) );
  nor2_1 U20904 ( .ip1(n21198), .ip2(n18535), .op(n18536) );
  nor2_1 U20905 ( .ip1(n18537), .ip2(n18536), .op(\pipeline/csr/N2099 ) );
  nand2_1 U20906 ( .ip1(\pipeline/csr/mscratch [18]), .ip2(n22013), .op(n18539) );
  nand2_1 U20907 ( .ip1(n22014), .ip2(n18563), .op(n18538) );
  nand2_1 U20908 ( .ip1(n18539), .ip2(n18538), .op(n9910) );
  nand2_1 U20909 ( .ip1(\pipeline/csr/from_host [18]), .ip2(n22372), .op(
        n18541) );
  nand2_1 U20910 ( .ip1(n22373), .ip2(n18563), .op(n18540) );
  nand2_1 U20911 ( .ip1(n18541), .ip2(n18540), .op(n9942) );
  nand2_1 U20912 ( .ip1(n22378), .ip2(n18563), .op(n18543) );
  nand2_1 U20913 ( .ip1(\pipeline/csr/to_host [18]), .ip2(n22376), .op(n18542)
         );
  nand2_1 U20914 ( .ip1(n18543), .ip2(n18542), .op(n8754) );
  or2_1 U20915 ( .ip1(n19804), .ip2(n21210), .op(n22244) );
  nor2_1 U20916 ( .ip1(n18572), .ip2(n22244), .op(n18546) );
  inv_1 U20917 ( .ip(\pipeline/csr/mtime_full [48]), .op(n19927) );
  inv_1 U20918 ( .ip(\pipeline/csr/mtime_full [46]), .op(n22174) );
  inv_1 U20919 ( .ip(\pipeline/csr/mtime_full [42]), .op(n19808) );
  nand2_1 U20920 ( .ip1(\pipeline/csr/mtime_full [41]), .ip2(n19722), .op(
        n19807) );
  nor2_1 U20921 ( .ip1(n19808), .ip2(n19807), .op(n22157) );
  nand2_1 U20922 ( .ip1(\pipeline/csr/mtime_full [43]), .ip2(n22157), .op(
        n22162) );
  nor2_1 U20923 ( .ip1(n22163), .ip2(n22162), .op(n22167) );
  nand2_1 U20924 ( .ip1(\pipeline/csr/mtime_full [45]), .ip2(n22167), .op(
        n22173) );
  nor2_1 U20925 ( .ip1(n22174), .ip2(n22173), .op(n22178) );
  nand2_1 U20926 ( .ip1(\pipeline/csr/mtime_full [47]), .ip2(n22178), .op(
        n22180) );
  nor2_1 U20927 ( .ip1(n19927), .ip2(n22180), .op(n22184) );
  nand2_1 U20928 ( .ip1(\pipeline/csr/mtime_full [49]), .ip2(n22184), .op(
        n22186) );
  inv_1 U20929 ( .ip(\pipeline/csr/mtime_full [50]), .op(n18544) );
  nor2_1 U20930 ( .ip1(n18544), .ip2(n22186), .op(n22190) );
  inv_1 U20931 ( .ip(n18449), .op(n22247) );
  not_ab_or_c_or_d U20932 ( .ip1(n22186), .ip2(n18544), .ip3(n22190), .ip4(
        n22247), .op(n18545) );
  or2_1 U20933 ( .ip1(n18546), .ip2(n18545), .op(\pipeline/csr/N2131 ) );
  inv_1 U20934 ( .ip(n21215), .op(n18547) );
  nor2_1 U20935 ( .ip1(n18547), .ip2(n21217), .op(n21145) );
  or2_1 U20936 ( .ip1(\pipeline/csr/cycle_full [18]), .ip2(n19988), .op(n18548) );
  nand2_1 U20937 ( .ip1(n18606), .ip2(n18548), .op(n18549) );
  or2_1 U20938 ( .ip1(n21145), .ip2(n18549), .op(n18551) );
  nor2_1 U20939 ( .ip1(n18605), .ip2(n21210), .op(n22021) );
  nand2_1 U20940 ( .ip1(n22021), .ip2(n18563), .op(n18550) );
  nand2_1 U20941 ( .ip1(n18551), .ip2(n18550), .op(\pipeline/csr/N1891 ) );
  nand2_1 U20942 ( .ip1(\pipeline/csr/mtimecmp [18]), .ip2(n22363), .op(n18553) );
  nand2_1 U20943 ( .ip1(n22365), .ip2(n18563), .op(n18552) );
  nand2_1 U20944 ( .ip1(n18553), .ip2(n18552), .op(n10004) );
  mux2_1 U20945 ( .ip1(\pipeline/csr/instret_full [18]), .ip2(n18558), .s(
        n18554), .op(n18557) );
  inv_1 U20946 ( .ip(n18555), .op(n21012) );
  nor2_1 U20947 ( .ip1(n21012), .ip2(n21011), .op(n18556) );
  nor2_1 U20948 ( .ip1(n18557), .ip2(n18556), .op(n18560) );
  nor2_1 U20949 ( .ip1(n18558), .ip2(n20990), .op(n18559) );
  nor2_1 U20950 ( .ip1(n18560), .ip2(n18559), .op(n18562) );
  nand2_1 U20951 ( .ip1(n21019), .ip2(n18563), .op(n18561) );
  nand2_1 U20952 ( .ip1(n18562), .ip2(n18561), .op(n10120) );
  nand2_1 U20953 ( .ip1(\pipeline/csr/mie [18]), .ip2(n22356), .op(n18565) );
  nand2_1 U20954 ( .ip1(n22357), .ip2(n18563), .op(n18564) );
  nand2_1 U20955 ( .ip1(n18565), .ip2(n18564), .op(n10042) );
  inv_1 U20956 ( .ip(\pipeline/csr/cycle_full [50]), .op(n18567) );
  nor2_1 U20957 ( .ip1(n19999), .ip2(n18567), .op(n18566) );
  not_ab_or_c_or_d U20958 ( .ip1(n19999), .ip2(n18567), .ip3(n18566), .ip4(
        n22314), .op(n18571) );
  nor2_1 U20959 ( .ip1(n18572), .ip2(n18568), .op(n18569) );
  inv_1 U20960 ( .ip(n22308), .op(n22316) );
  nor2_1 U20961 ( .ip1(n18569), .ip2(n22316), .op(n18570) );
  nor2_1 U20962 ( .ip1(n18571), .ip2(n18570), .op(\pipeline/csr/N1923 ) );
  nor2_1 U20963 ( .ip1(n18572), .ip2(n21110), .op(n18576) );
  inv_1 U20964 ( .ip(\pipeline/csr/instret_full [50]), .op(n18574) );
  nor2_1 U20965 ( .ip1(n18574), .ip2(n18573), .op(n18626) );
  not_ab_or_c_or_d U20966 ( .ip1(n18574), .ip2(n18573), .ip3(n21111), .ip4(
        n18626), .op(n18575) );
  ab_or_c_or_d U20967 ( .ip1(n21117), .ip2(\pipeline/csr/instret_full [50]), 
        .ip3(n18576), .ip4(n18575), .op(n10088) );
  nand2_1 U20968 ( .ip1(n21032), .ip2(n22189), .op(n18578) );
  nand2_1 U20969 ( .ip1(\pipeline/csr/mtvec [19]), .ip2(n20705), .op(n18577)
         );
  nand2_1 U20970 ( .ip1(n18578), .ip2(n18577), .op(n9973) );
  mux2_1 U20971 ( .ip1(\pipeline/PC_WB [19]), .ip2(\pipeline/PC_DX [19]), .s(
        n17777), .op(n8884) );
  nand2_1 U20972 ( .ip1(dmem_rdata[19]), .ip2(n21585), .op(n18582) );
  nand2_1 U20973 ( .ip1(n18579), .ip2(n21583), .op(n18581) );
  nand2_1 U20974 ( .ip1(dmem_rdata[27]), .ip2(n19324), .op(n18580) );
  nand4_1 U20975 ( .ip1(n21588), .ip2(n18582), .ip3(n18581), .ip4(n18580), 
        .op(n18583) );
  mux2_1 U20976 ( .ip1(\pipeline/regfile/data[29][19] ), .ip2(n18583), .s(
        n21619), .op(n8981) );
  mux2_1 U20977 ( .ip1(\pipeline/regfile/data[14][19] ), .ip2(n18583), .s(
        n21604), .op(n9461) );
  mux2_1 U20978 ( .ip1(\pipeline/regfile/data[22][19] ), .ip2(n18583), .s(
        n21589), .op(n9205) );
  mux2_1 U20979 ( .ip1(\pipeline/regfile/data[5][19] ), .ip2(n18583), .s(
        n21598), .op(n9749) );
  mux2_1 U20980 ( .ip1(\pipeline/regfile/data[27][19] ), .ip2(n18583), .s(
        n21612), .op(n9045) );
  mux2_1 U20981 ( .ip1(\pipeline/regfile/data[26][19] ), .ip2(n18583), .s(
        n21607), .op(n9077) );
  mux2_1 U20982 ( .ip1(\pipeline/regfile/data[28][19] ), .ip2(n18583), .s(
        n21590), .op(n9013) );
  mux2_1 U20983 ( .ip1(\pipeline/regfile/data[31][19] ), .ip2(n18583), .s(
        n21606), .op(n8917) );
  mux2_1 U20984 ( .ip1(\pipeline/regfile/data[19][19] ), .ip2(n18583), .s(
        n21592), .op(n9301) );
  mux2_1 U20985 ( .ip1(\pipeline/regfile/data[6][19] ), .ip2(n18583), .s(
        n21597), .op(n9717) );
  mux2_1 U20986 ( .ip1(\pipeline/regfile/data[30][19] ), .ip2(n18583), .s(
        n21594), .op(n8949) );
  mux2_1 U20987 ( .ip1(\pipeline/regfile/data[18][19] ), .ip2(n18583), .s(
        n21595), .op(n9333) );
  mux2_1 U20988 ( .ip1(\pipeline/regfile/data[11][19] ), .ip2(n18583), .s(
        n21593), .op(n9557) );
  mux2_1 U20989 ( .ip1(\pipeline/regfile/data[25][19] ), .ip2(n18583), .s(
        n21602), .op(n9109) );
  mux2_1 U20990 ( .ip1(\pipeline/regfile/data[13][19] ), .ip2(n18583), .s(
        n21600), .op(n9493) );
  mux2_1 U20991 ( .ip1(\pipeline/regfile/data[17][19] ), .ip2(n18583), .s(
        n21616), .op(n9365) );
  mux2_1 U20992 ( .ip1(\pipeline/regfile/data[23][19] ), .ip2(n18583), .s(
        n21596), .op(n9173) );
  mux2_1 U20993 ( .ip1(\pipeline/regfile/data[12][19] ), .ip2(n18583), .s(
        n21591), .op(n9525) );
  mux2_1 U20994 ( .ip1(\pipeline/regfile/data[7][19] ), .ip2(n18583), .s(
        n21614), .op(n9685) );
  mux2_1 U20995 ( .ip1(\pipeline/regfile/data[8][19] ), .ip2(n18583), .s(
        n21617), .op(n9653) );
  mux2_1 U20996 ( .ip1(\pipeline/regfile/data[15][19] ), .ip2(n18583), .s(
        n21613), .op(n9429) );
  mux2_1 U20997 ( .ip1(\pipeline/regfile/data[10][19] ), .ip2(n18583), .s(
        n21618), .op(n9589) );
  mux2_1 U20998 ( .ip1(\pipeline/regfile/data[21][19] ), .ip2(n18583), .s(
        n21615), .op(n9237) );
  mux2_1 U20999 ( .ip1(\pipeline/regfile/data[24][19] ), .ip2(n18583), .s(
        n21603), .op(n9141) );
  mux2_1 U21000 ( .ip1(\pipeline/regfile/data[20][19] ), .ip2(n18583), .s(
        n21601), .op(n9269) );
  mux2_1 U21001 ( .ip1(\pipeline/regfile/data[9][19] ), .ip2(n18583), .s(
        n21609), .op(n9621) );
  mux2_1 U21002 ( .ip1(\pipeline/regfile/data[16][19] ), .ip2(n18583), .s(
        n21608), .op(n9397) );
  mux2_1 U21003 ( .ip1(\pipeline/regfile/data[3][19] ), .ip2(n18583), .s(
        n21599), .op(n9813) );
  mux2_1 U21004 ( .ip1(\pipeline/regfile/data[1][19] ), .ip2(n18583), .s(
        n21611), .op(n9877) );
  mux2_1 U21005 ( .ip1(\pipeline/regfile/data[2][19] ), .ip2(n18583), .s(
        n21610), .op(n9845) );
  mux2_1 U21006 ( .ip1(\pipeline/regfile/data[4][19] ), .ip2(n18583), .s(
        n21605), .op(n9781) );
  mux2_1 U21007 ( .ip1(dmem_haddr[19]), .ip2(\pipeline/alu_out_WB [19]), .s(
        n19505), .op(n8713) );
  inv_1 U21008 ( .ip(n22189), .op(n20027) );
  nor2_1 U21009 ( .ip1(n20027), .ip2(n22267), .op(n18587) );
  not_ab_or_c_or_d U21010 ( .ip1(n18585), .ip2(n18584), .ip3(n19508), .ip4(
        n22276), .op(n18586) );
  or2_1 U21011 ( .ip1(n18587), .ip2(n18586), .op(\pipeline/csr/N1988 ) );
  inv_1 U21012 ( .ip(n18588), .op(n18589) );
  nor2_1 U21013 ( .ip1(\pipeline/csr/time_full [19]), .ip2(n18589), .op(n18591) );
  nor3_1 U21014 ( .ip1(n21177), .ip2(n19512), .ip3(n18591), .op(n18590) );
  not_ab_or_c_or_d U21015 ( .ip1(n21179), .ip2(n22189), .ip3(n21217), .ip4(
        n18590), .op(n18594) );
  nor2_1 U21016 ( .ip1(n18591), .ip2(n19512), .op(n18592) );
  nor2_1 U21017 ( .ip1(n22254), .ip2(n18592), .op(n18593) );
  nor2_1 U21018 ( .ip1(n18594), .ip2(n18593), .op(\pipeline/csr/N1956 ) );
  nand2_1 U21019 ( .ip1(n22008), .ip2(n22189), .op(n18598) );
  xor2_1 U21020 ( .ip1(n18595), .ip2(\pipeline/csr/mtime_full [19]), .op(
        n18596) );
  nand2_1 U21021 ( .ip1(n18596), .ip2(n22009), .op(n18597) );
  nand2_1 U21022 ( .ip1(n18598), .ip2(n18597), .op(\pipeline/csr/N2100 ) );
  nand2_1 U21023 ( .ip1(\pipeline/csr/mscratch [19]), .ip2(n22013), .op(n18600) );
  nand2_1 U21024 ( .ip1(n22014), .ip2(n22189), .op(n18599) );
  nand2_1 U21025 ( .ip1(n18600), .ip2(n18599), .op(n9909) );
  nand2_1 U21026 ( .ip1(\pipeline/csr/from_host [19]), .ip2(n22372), .op(
        n18602) );
  nand2_1 U21027 ( .ip1(n22373), .ip2(n22189), .op(n18601) );
  nand2_1 U21028 ( .ip1(n18602), .ip2(n18601), .op(n9941) );
  nand2_1 U21029 ( .ip1(n22378), .ip2(n22189), .op(n18604) );
  nand2_1 U21030 ( .ip1(\pipeline/csr/to_host [19]), .ip2(n22376), .op(n18603)
         );
  nand2_1 U21031 ( .ip1(n18604), .ip2(n18603), .op(n8753) );
  inv_1 U21032 ( .ip(n18605), .op(n21076) );
  inv_1 U21033 ( .ip(n18606), .op(n18607) );
  nor2_1 U21034 ( .ip1(\pipeline/csr/cycle_full [19]), .ip2(n18607), .op(
        n18609) );
  nor3_1 U21035 ( .ip1(n19532), .ip2(n18609), .ip3(n21215), .op(n18608) );
  not_ab_or_c_or_d U21036 ( .ip1(n21076), .ip2(n22189), .ip3(n21217), .ip4(
        n18608), .op(n18612) );
  nor2_1 U21037 ( .ip1(n18609), .ip2(n19532), .op(n18610) );
  nor2_1 U21038 ( .ip1(n21198), .ip2(n18610), .op(n18611) );
  nor2_1 U21039 ( .ip1(n18612), .ip2(n18611), .op(\pipeline/csr/N1892 ) );
  nand2_1 U21040 ( .ip1(\pipeline/csr/mtimecmp [19]), .ip2(n22363), .op(n18614) );
  nand2_1 U21041 ( .ip1(n22365), .ip2(n22189), .op(n18613) );
  nand2_1 U21042 ( .ip1(n18614), .ip2(n18613), .op(n10003) );
  nor2_1 U21043 ( .ip1(n20027), .ip2(n21001), .op(n18619) );
  inv_1 U21044 ( .ip(\pipeline/csr/instret_full [19]), .op(n18616) );
  mux2_1 U21045 ( .ip1(n18616), .ip2(\pipeline/csr/instret_full [19]), .s(
        n18615), .op(n18617) );
  nor2_1 U21046 ( .ip1(n21005), .ip2(n18617), .op(n18618) );
  ab_or_c_or_d U21047 ( .ip1(n21016), .ip2(\pipeline/csr/instret_full [19]), 
        .ip3(n18619), .ip4(n18618), .op(n10119) );
  nand2_1 U21048 ( .ip1(\pipeline/csr/mie [19]), .ip2(n22356), .op(n18621) );
  nand2_1 U21049 ( .ip1(n22357), .ip2(n22189), .op(n18620) );
  nand2_1 U21050 ( .ip1(n18621), .ip2(n18620), .op(n10041) );
  nor2_1 U21051 ( .ip1(n20027), .ip2(n22305), .op(n18625) );
  not_ab_or_c_or_d U21052 ( .ip1(n18623), .ip2(n18622), .ip3(n19550), .ip4(
        n22308), .op(n18624) );
  or2_1 U21053 ( .ip1(n18625), .ip2(n18624), .op(\pipeline/csr/N1924 ) );
  nand2_1 U21054 ( .ip1(n20844), .ip2(n22189), .op(n18630) );
  nand2_1 U21055 ( .ip1(\pipeline/csr/instret_full [51]), .ip2(n21117), .op(
        n18629) );
  nand2_1 U21056 ( .ip1(\pipeline/csr/instret_full [51]), .ip2(n18626), .op(
        n18631) );
  or2_1 U21057 ( .ip1(\pipeline/csr/instret_full [51]), .ip2(n18626), .op(
        n18627) );
  nand3_1 U21058 ( .ip1(n18631), .ip2(n20334), .ip3(n18627), .op(n18628) );
  nand3_1 U21059 ( .ip1(n18630), .ip2(n18629), .ip3(n18628), .op(n10087) );
  nand2_1 U21060 ( .ip1(n19549), .ip2(n20844), .op(n18636) );
  and2_1 U21061 ( .ip1(n21117), .ip2(\pipeline/csr/instret_full [52]), .op(
        n18634) );
  inv_1 U21062 ( .ip(\pipeline/csr/instret_full [52]), .op(n18632) );
  nor2_1 U21063 ( .ip1(n18632), .ip2(n18631), .op(n18700) );
  not_ab_or_c_or_d U21064 ( .ip1(n18632), .ip2(n18631), .ip3(n18700), .ip4(
        n21111), .op(n18633) );
  nor2_1 U21065 ( .ip1(n18634), .ip2(n18633), .op(n18635) );
  nand2_1 U21066 ( .ip1(n18636), .ip2(n18635), .op(n10086) );
  nor2_1 U21067 ( .ip1(n18638), .ip2(n18637), .op(n18641) );
  xor2_1 U21068 ( .ip1(\pipeline/PC_WB [21]), .ip2(n20051), .op(n18639) );
  nor2_1 U21069 ( .ip1(n21171), .ip2(n18639), .op(n18640) );
  ab_or_c_or_d U21070 ( .ip1(n21043), .ip2(n22368), .ip3(n18641), .ip4(n18640), 
        .op(n8850) );
  nor2_1 U21071 ( .ip1(n22368), .ip2(n21029), .op(n18645) );
  inv_1 U21072 ( .ip(\pipeline/csr/mtvec [21]), .op(n18642) );
  nor2_1 U21073 ( .ip1(n21089), .ip2(n18642), .op(n18643) );
  nor2_1 U21074 ( .ip1(n21032), .ip2(n18643), .op(n18644) );
  nor2_1 U21075 ( .ip1(n18645), .ip2(n18644), .op(n9971) );
  nand2_1 U21076 ( .ip1(dmem_rdata[21]), .ip2(n21585), .op(n18649) );
  nand2_1 U21077 ( .ip1(n18646), .ip2(n21583), .op(n18648) );
  nand2_1 U21078 ( .ip1(dmem_rdata[29]), .ip2(n19324), .op(n18647) );
  nand4_1 U21079 ( .ip1(n21588), .ip2(n18649), .ip3(n18648), .ip4(n18647), 
        .op(n18650) );
  mux2_1 U21080 ( .ip1(\pipeline/regfile/data[29][21] ), .ip2(n18650), .s(
        n19353), .op(n8979) );
  mux2_1 U21081 ( .ip1(\pipeline/regfile/data[14][21] ), .ip2(n18650), .s(
        n19354), .op(n9459) );
  mux2_1 U21082 ( .ip1(\pipeline/regfile/data[22][21] ), .ip2(n18650), .s(
        n19355), .op(n9203) );
  mux2_1 U21083 ( .ip1(\pipeline/regfile/data[5][21] ), .ip2(n18650), .s(
        n19356), .op(n9747) );
  mux2_1 U21084 ( .ip1(\pipeline/regfile/data[27][21] ), .ip2(n18650), .s(
        n19357), .op(n9043) );
  mux2_1 U21085 ( .ip1(\pipeline/regfile/data[26][21] ), .ip2(n18650), .s(
        n19358), .op(n9075) );
  mux2_1 U21086 ( .ip1(\pipeline/regfile/data[28][21] ), .ip2(n18650), .s(
        n19359), .op(n9011) );
  mux2_1 U21087 ( .ip1(\pipeline/regfile/data[31][21] ), .ip2(n18650), .s(
        n19360), .op(n8915) );
  mux2_1 U21088 ( .ip1(\pipeline/regfile/data[19][21] ), .ip2(n18650), .s(
        n19361), .op(n9299) );
  mux2_1 U21089 ( .ip1(\pipeline/regfile/data[6][21] ), .ip2(n18650), .s(
        n19362), .op(n9715) );
  mux2_1 U21090 ( .ip1(\pipeline/regfile/data[30][21] ), .ip2(n18650), .s(
        n19363), .op(n8947) );
  mux2_1 U21091 ( .ip1(\pipeline/regfile/data[18][21] ), .ip2(n18650), .s(
        n19364), .op(n9331) );
  mux2_1 U21092 ( .ip1(\pipeline/regfile/data[11][21] ), .ip2(n18650), .s(
        n19365), .op(n9555) );
  mux2_1 U21093 ( .ip1(\pipeline/regfile/data[25][21] ), .ip2(n18650), .s(
        n19366), .op(n9107) );
  mux2_1 U21094 ( .ip1(\pipeline/regfile/data[13][21] ), .ip2(n18650), .s(
        n19367), .op(n9491) );
  mux2_1 U21095 ( .ip1(\pipeline/regfile/data[17][21] ), .ip2(n18650), .s(
        n19368), .op(n9363) );
  mux2_1 U21096 ( .ip1(\pipeline/regfile/data[23][21] ), .ip2(n18650), .s(
        n19369), .op(n9171) );
  mux2_1 U21097 ( .ip1(\pipeline/regfile/data[12][21] ), .ip2(n18650), .s(
        n19370), .op(n9523) );
  mux2_1 U21098 ( .ip1(\pipeline/regfile/data[7][21] ), .ip2(n18650), .s(
        n19371), .op(n9683) );
  mux2_1 U21099 ( .ip1(\pipeline/regfile/data[8][21] ), .ip2(n18650), .s(
        n19372), .op(n9651) );
  mux2_1 U21100 ( .ip1(\pipeline/regfile/data[15][21] ), .ip2(n18650), .s(
        n19373), .op(n9427) );
  mux2_1 U21101 ( .ip1(\pipeline/regfile/data[10][21] ), .ip2(n18650), .s(
        n19374), .op(n9587) );
  mux2_1 U21102 ( .ip1(\pipeline/regfile/data[21][21] ), .ip2(n18650), .s(
        n19375), .op(n9235) );
  mux2_1 U21103 ( .ip1(\pipeline/regfile/data[24][21] ), .ip2(n18650), .s(
        n19376), .op(n9139) );
  mux2_1 U21104 ( .ip1(\pipeline/regfile/data[20][21] ), .ip2(n18650), .s(
        n19377), .op(n9267) );
  mux2_1 U21105 ( .ip1(\pipeline/regfile/data[9][21] ), .ip2(n18650), .s(
        n19378), .op(n9619) );
  mux2_1 U21106 ( .ip1(\pipeline/regfile/data[16][21] ), .ip2(n18650), .s(
        n19379), .op(n9395) );
  mux2_1 U21107 ( .ip1(\pipeline/regfile/data[3][21] ), .ip2(n18650), .s(
        n19380), .op(n9811) );
  mux2_1 U21108 ( .ip1(\pipeline/regfile/data[1][21] ), .ip2(n18650), .s(
        n19381), .op(n9875) );
  mux2_1 U21109 ( .ip1(\pipeline/regfile/data[2][21] ), .ip2(n18650), .s(
        n19382), .op(n9843) );
  mux2_1 U21110 ( .ip1(\pipeline/regfile/data[4][21] ), .ip2(n18650), .s(
        n19383), .op(n9779) );
  mux2_1 U21111 ( .ip1(dmem_haddr[21]), .ip2(\pipeline/alu_out_WB [21]), .s(
        n19505), .op(n8711) );
  nand2_1 U21112 ( .ip1(n22282), .ip2(n22368), .op(n18654) );
  xnor2_1 U21113 ( .ip1(\pipeline/csr/time_full [53]), .ip2(n18651), .op(
        n18652) );
  nand2_1 U21114 ( .ip1(n22284), .ip2(n18652), .op(n18653) );
  nand2_1 U21115 ( .ip1(n18654), .ip2(n18653), .op(\pipeline/csr/N1990 ) );
  inv_1 U21116 ( .ip(n18655), .op(n18656) );
  nor2_1 U21117 ( .ip1(\pipeline/csr/time_full [21]), .ip2(n18656), .op(n18658) );
  nor3_1 U21118 ( .ip1(n21177), .ip2(n20063), .ip3(n18658), .op(n18657) );
  not_ab_or_c_or_d U21119 ( .ip1(n21179), .ip2(n22368), .ip3(n21217), .ip4(
        n18657), .op(n18661) );
  nor2_1 U21120 ( .ip1(n18658), .ip2(n20063), .op(n18659) );
  nor2_1 U21121 ( .ip1(n21198), .ip2(n18659), .op(n18660) );
  nor2_1 U21122 ( .ip1(n18661), .ip2(n18660), .op(\pipeline/csr/N1958 ) );
  inv_1 U21123 ( .ip(\pipeline/csr/mtime_full [21]), .op(n19661) );
  xor2_1 U21124 ( .ip1(n19521), .ip2(n19661), .op(n18663) );
  nor2_1 U21125 ( .ip1(n21193), .ip2(n18663), .op(n18662) );
  not_ab_or_c_or_d U21126 ( .ip1(n21195), .ip2(n22368), .ip3(n21217), .ip4(
        n18662), .op(n18666) );
  inv_1 U21127 ( .ip(n18663), .op(n18664) );
  nor2_1 U21128 ( .ip1(n21198), .ip2(n18664), .op(n18665) );
  nor2_1 U21129 ( .ip1(n18666), .ip2(n18665), .op(\pipeline/csr/N2102 ) );
  nand2_1 U21130 ( .ip1(\pipeline/csr/mscratch [21]), .ip2(n22013), .op(n18668) );
  nand2_1 U21131 ( .ip1(n22014), .ip2(n22368), .op(n18667) );
  nand2_1 U21132 ( .ip1(n18668), .ip2(n18667), .op(n9907) );
  nand2_1 U21133 ( .ip1(\pipeline/csr/from_host [21]), .ip2(n22372), .op(
        n18670) );
  nand2_1 U21134 ( .ip1(n22373), .ip2(n22368), .op(n18669) );
  nand2_1 U21135 ( .ip1(n18670), .ip2(n18669), .op(n9939) );
  nand2_1 U21136 ( .ip1(n22378), .ip2(n22368), .op(n18672) );
  nand2_1 U21137 ( .ip1(\pipeline/csr/to_host [21]), .ip2(n22376), .op(n18671)
         );
  nand2_1 U21138 ( .ip1(n18672), .ip2(n18671), .op(n8751) );
  inv_1 U21139 ( .ip(n19534), .op(n18673) );
  nor2_1 U21140 ( .ip1(\pipeline/csr/cycle_full [21]), .ip2(n18673), .op(
        n18675) );
  nor3_1 U21141 ( .ip1(n20083), .ip2(n18675), .ip3(n21215), .op(n18674) );
  not_ab_or_c_or_d U21142 ( .ip1(n21076), .ip2(n22368), .ip3(n21217), .ip4(
        n18674), .op(n18678) );
  nor2_1 U21143 ( .ip1(n18675), .ip2(n20083), .op(n18676) );
  nor2_1 U21144 ( .ip1(n21198), .ip2(n18676), .op(n18677) );
  nor2_1 U21145 ( .ip1(n18678), .ip2(n18677), .op(\pipeline/csr/N1894 ) );
  inv_1 U21146 ( .ip(\pipeline/csr/instret_full [21]), .op(n18680) );
  nor2_1 U21147 ( .ip1(n18680), .ip2(n20990), .op(n18683) );
  mux2_1 U21148 ( .ip1(n18680), .ip2(\pipeline/csr/instret_full [21]), .s(
        n18679), .op(n18681) );
  nor2_1 U21149 ( .ip1(n21005), .ip2(n18681), .op(n18682) );
  ab_or_c_or_d U21150 ( .ip1(n21019), .ip2(n22368), .ip3(n18683), .ip4(n18682), 
        .op(n10117) );
  nand2_1 U21151 ( .ip1(\pipeline/csr/mie [21]), .ip2(n22356), .op(n18685) );
  nand2_1 U21152 ( .ip1(n22357), .ip2(n22368), .op(n18684) );
  nand2_1 U21153 ( .ip1(n18685), .ip2(n18684), .op(n10039) );
  inv_1 U21154 ( .ip(n22368), .op(n18686) );
  inv_1 U21155 ( .ip(n22314), .op(n22305) );
  nor2_1 U21156 ( .ip1(n18686), .ip2(n22305), .op(n18689) );
  not_ab_or_c_or_d U21157 ( .ip1(n19552), .ip2(n18687), .ip3(n20101), .ip4(
        n22308), .op(n18688) );
  or2_1 U21158 ( .ip1(n18689), .ip2(n18688), .op(\pipeline/csr/N1926 ) );
  xor2_1 U21159 ( .ip1(\pipeline/csr/instret_full [53]), .ip2(n18700), .op(
        n18696) );
  nand2_1 U21160 ( .ip1(n18696), .ip2(n18690), .op(n18693) );
  nand2_1 U21161 ( .ip1(n18691), .ip2(n22368), .op(n18692) );
  nand2_1 U21162 ( .ip1(n18693), .ip2(n18692), .op(n18694) );
  nand2_1 U21163 ( .ip1(n18695), .ip2(n18694), .op(n18699) );
  nand2_1 U21164 ( .ip1(\pipeline/csr/instret_full [53]), .ip2(n21117), .op(
        n18698) );
  nand2_1 U21165 ( .ip1(n18696), .ip2(n21011), .op(n18697) );
  nand3_1 U21166 ( .ip1(n18699), .ip2(n18698), .ip3(n18697), .op(n10085) );
  inv_1 U21167 ( .ip(n20100), .op(n22203) );
  nor2_1 U21168 ( .ip1(n22203), .ip2(n21110), .op(n18704) );
  inv_1 U21169 ( .ip(\pipeline/csr/instret_full [54]), .op(n18702) );
  nand2_1 U21170 ( .ip1(n18700), .ip2(\pipeline/csr/instret_full [53]), .op(
        n18701) );
  and3_1 U21171 ( .ip1(n18700), .ip2(\pipeline/csr/instret_full [53]), .ip3(
        \pipeline/csr/instret_full [54]), .op(n18705) );
  not_ab_or_c_or_d U21172 ( .ip1(n18702), .ip2(n18701), .ip3(n18705), .ip4(
        n21111), .op(n18703) );
  ab_or_c_or_d U21173 ( .ip1(\pipeline/csr/instret_full [54]), .ip2(n21117), 
        .ip3(n18704), .ip4(n18703), .op(n10084) );
  nand2_1 U21174 ( .ip1(n20844), .ip2(n22274), .op(n18709) );
  nand2_1 U21175 ( .ip1(n21117), .ip2(\pipeline/csr/instret_full [55]), .op(
        n18708) );
  nand2_1 U21176 ( .ip1(\pipeline/csr/instret_full [55]), .ip2(n18705), .op(
        n18798) );
  or2_1 U21177 ( .ip1(\pipeline/csr/instret_full [55]), .ip2(n18705), .op(
        n18706) );
  nand3_1 U21178 ( .ip1(n20334), .ip2(n18798), .ip3(n18706), .op(n18707) );
  nand3_1 U21179 ( .ip1(n18709), .ip2(n18708), .ip3(n18707), .op(n10083) );
  inv_1 U21180 ( .ip(n18794), .op(n22212) );
  nor2_1 U21181 ( .ip1(n22212), .ip2(n21168), .op(n18712) );
  xor2_1 U21182 ( .ip1(\pipeline/PC_WB [24]), .ip2(n18827), .op(n18710) );
  nor2_1 U21183 ( .ip1(n21171), .ip2(n18710), .op(n18711) );
  ab_or_c_or_d U21184 ( .ip1(n21174), .ip2(\pipeline/epc [24]), .ip3(n18712), 
        .ip4(n18711), .op(n8847) );
  nor2_1 U21185 ( .ip1(n18794), .ip2(n21029), .op(n18716) );
  inv_1 U21186 ( .ip(\pipeline/csr/mtvec [24]), .op(n18713) );
  nor2_1 U21187 ( .ip1(n21089), .ip2(n18713), .op(n18714) );
  nor2_1 U21188 ( .ip1(n21032), .ip2(n18714), .op(n18715) );
  nor2_1 U21189 ( .ip1(n18716), .ip2(n18715), .op(n9968) );
  nand2_1 U21190 ( .ip1(n18717), .ip2(n21583), .op(n18719) );
  nand2_1 U21191 ( .ip1(n21585), .ip2(dmem_rdata[24]), .op(n18718) );
  nand3_1 U21192 ( .ip1(n21588), .ip2(n18719), .ip3(n18718), .op(n18720) );
  mux2_1 U21193 ( .ip1(\pipeline/regfile/data[29][24] ), .ip2(n18720), .s(
        n19353), .op(n8976) );
  mux2_1 U21194 ( .ip1(\pipeline/regfile/data[14][24] ), .ip2(n18720), .s(
        n19354), .op(n9456) );
  mux2_1 U21195 ( .ip1(\pipeline/regfile/data[22][24] ), .ip2(n18720), .s(
        n19355), .op(n9200) );
  mux2_1 U21196 ( .ip1(\pipeline/regfile/data[5][24] ), .ip2(n18720), .s(
        n19356), .op(n9744) );
  mux2_1 U21197 ( .ip1(\pipeline/regfile/data[27][24] ), .ip2(n18720), .s(
        n19357), .op(n9040) );
  mux2_1 U21198 ( .ip1(\pipeline/regfile/data[26][24] ), .ip2(n18720), .s(
        n19358), .op(n9072) );
  mux2_1 U21199 ( .ip1(\pipeline/regfile/data[28][24] ), .ip2(n18720), .s(
        n19359), .op(n9008) );
  mux2_1 U21200 ( .ip1(\pipeline/regfile/data[31][24] ), .ip2(n18720), .s(
        n19360), .op(n8912) );
  mux2_1 U21201 ( .ip1(\pipeline/regfile/data[19][24] ), .ip2(n18720), .s(
        n19361), .op(n9296) );
  mux2_1 U21202 ( .ip1(\pipeline/regfile/data[6][24] ), .ip2(n18720), .s(
        n19362), .op(n9712) );
  mux2_1 U21203 ( .ip1(\pipeline/regfile/data[30][24] ), .ip2(n18720), .s(
        n19363), .op(n8944) );
  mux2_1 U21204 ( .ip1(\pipeline/regfile/data[18][24] ), .ip2(n18720), .s(
        n19364), .op(n9328) );
  mux2_1 U21205 ( .ip1(\pipeline/regfile/data[11][24] ), .ip2(n18720), .s(
        n19365), .op(n9552) );
  mux2_1 U21206 ( .ip1(\pipeline/regfile/data[25][24] ), .ip2(n18720), .s(
        n19366), .op(n9104) );
  mux2_1 U21207 ( .ip1(\pipeline/regfile/data[13][24] ), .ip2(n18720), .s(
        n19367), .op(n9488) );
  mux2_1 U21208 ( .ip1(\pipeline/regfile/data[17][24] ), .ip2(n18720), .s(
        n19368), .op(n9360) );
  mux2_1 U21209 ( .ip1(\pipeline/regfile/data[23][24] ), .ip2(n18720), .s(
        n19369), .op(n9168) );
  mux2_1 U21210 ( .ip1(\pipeline/regfile/data[12][24] ), .ip2(n18720), .s(
        n19370), .op(n9520) );
  mux2_1 U21211 ( .ip1(\pipeline/regfile/data[7][24] ), .ip2(n18720), .s(
        n19371), .op(n9680) );
  mux2_1 U21212 ( .ip1(\pipeline/regfile/data[8][24] ), .ip2(n18720), .s(
        n19372), .op(n9648) );
  mux2_1 U21213 ( .ip1(\pipeline/regfile/data[15][24] ), .ip2(n18720), .s(
        n19373), .op(n9424) );
  mux2_1 U21214 ( .ip1(\pipeline/regfile/data[10][24] ), .ip2(n18720), .s(
        n19374), .op(n9584) );
  mux2_1 U21215 ( .ip1(\pipeline/regfile/data[21][24] ), .ip2(n18720), .s(
        n19375), .op(n9232) );
  mux2_1 U21216 ( .ip1(\pipeline/regfile/data[24][24] ), .ip2(n18720), .s(
        n19376), .op(n9136) );
  mux2_1 U21217 ( .ip1(\pipeline/regfile/data[20][24] ), .ip2(n18720), .s(
        n19377), .op(n9264) );
  mux2_1 U21218 ( .ip1(\pipeline/regfile/data[9][24] ), .ip2(n18720), .s(
        n19378), .op(n9616) );
  mux2_1 U21219 ( .ip1(\pipeline/regfile/data[16][24] ), .ip2(n18720), .s(
        n19379), .op(n9392) );
  mux2_1 U21220 ( .ip1(\pipeline/regfile/data[3][24] ), .ip2(n18720), .s(
        n19380), .op(n9808) );
  mux2_1 U21221 ( .ip1(\pipeline/regfile/data[1][24] ), .ip2(n18720), .s(
        n19381), .op(n9872) );
  mux2_1 U21222 ( .ip1(\pipeline/regfile/data[2][24] ), .ip2(n18720), .s(
        n19382), .op(n9840) );
  mux2_1 U21223 ( .ip1(\pipeline/regfile/data[4][24] ), .ip2(n18720), .s(
        n19383), .op(n9776) );
  nand2_1 U21224 ( .ip1(n18722), .ip2(n18721), .op(n18727) );
  nand2_1 U21225 ( .ip1(n20878), .ip2(n18723), .op(n18724) );
  nand2_1 U21226 ( .ip1(n18725), .ip2(n18724), .op(n18726) );
  xnor2_1 U21227 ( .ip1(n18727), .ip2(n18726), .op(n18752) );
  nor2_1 U21228 ( .ip1(n20883), .ip2(n18728), .op(n18751) );
  nand2_1 U21229 ( .ip1(n18729), .ip2(n20736), .op(n18749) );
  nor3_1 U21230 ( .ip1(n18730), .ip2(n21551), .ip3(n13656), .op(n18734) );
  nor2_1 U21231 ( .ip1(n18731), .ip2(n10186), .op(n18732) );
  nor2_1 U21232 ( .ip1(n20907), .ip2(n18732), .op(n18733) );
  not_ab_or_c_or_d U21233 ( .ip1(n20911), .ip2(n18735), .ip3(n18734), .ip4(
        n18733), .op(n18747) );
  nor2_1 U21234 ( .ip1(n20885), .ip2(n19046), .op(n18736) );
  not_ab_or_c_or_d U21235 ( .ip1(n20896), .ip2(n19060), .ip3(n20724), .ip4(
        n18736), .op(n18745) );
  nand2_1 U21236 ( .ip1(n19059), .ip2(n21540), .op(n18744) );
  nand2_1 U21237 ( .ip1(n21536), .ip2(n18737), .op(n18742) );
  nand2_1 U21238 ( .ip1(n18927), .ip2(n10186), .op(n18741) );
  nand2_1 U21239 ( .ip1(n20892), .ip2(n18738), .op(n18740) );
  nand2_1 U21240 ( .ip1(n19056), .ip2(n17530), .op(n18739) );
  and4_1 U21241 ( .ip1(n18742), .ip2(n18741), .ip3(n18740), .ip4(n18739), .op(
        n19058) );
  nand2_1 U21242 ( .ip1(n19058), .ip2(n19427), .op(n18743) );
  nand3_1 U21243 ( .ip1(n18745), .ip2(n18744), .ip3(n18743), .op(n18746) );
  nand4_1 U21244 ( .ip1(n18749), .ip2(n18748), .ip3(n18747), .ip4(n18746), 
        .op(n18750) );
  ab_or_c_or_d U21245 ( .ip1(n18752), .ip2(n21577), .ip3(n18751), .ip4(n18750), 
        .op(dmem_haddr[24]) );
  mux2_1 U21246 ( .ip1(dmem_haddr[24]), .ip2(\pipeline/alu_out_WB [24]), .s(
        n19505), .op(n8708) );
  nand2_1 U21247 ( .ip1(n22282), .ip2(n18794), .op(n18755) );
  or2_1 U21248 ( .ip1(\pipeline/csr/time_full [56]), .ip2(n22275), .op(n18753)
         );
  nand3_1 U21249 ( .ip1(n18824), .ip2(n18753), .ip3(n22284), .op(n18754) );
  nand2_1 U21250 ( .ip1(n18755), .ip2(n18754), .op(\pipeline/csr/N1993 ) );
  or2_1 U21251 ( .ip1(\pipeline/csr/time_full [24]), .ip2(n20118), .op(n18756)
         );
  nand2_1 U21252 ( .ip1(n18757), .ip2(n18756), .op(n18758) );
  or2_1 U21253 ( .ip1(n22002), .ip2(n18758), .op(n18760) );
  nand2_1 U21254 ( .ip1(n22005), .ip2(n18794), .op(n18759) );
  nand2_1 U21255 ( .ip1(n18760), .ip2(n18759), .op(\pipeline/csr/N1961 ) );
  inv_1 U21256 ( .ip(n18761), .op(n18762) );
  nor2_1 U21257 ( .ip1(\pipeline/csr/mtime_full [24]), .ip2(n18762), .op(
        n18764) );
  nor3_1 U21258 ( .ip1(n21193), .ip2(n18764), .ip3(n18807), .op(n18763) );
  not_ab_or_c_or_d U21259 ( .ip1(n21195), .ip2(n18794), .ip3(n21217), .ip4(
        n18763), .op(n18767) );
  nor2_1 U21260 ( .ip1(n18764), .ip2(n18807), .op(n18765) );
  nor2_1 U21261 ( .ip1(n21198), .ip2(n18765), .op(n18766) );
  nor2_1 U21262 ( .ip1(n18767), .ip2(n18766), .op(\pipeline/csr/N2105 ) );
  nand2_1 U21263 ( .ip1(\pipeline/csr/mscratch [24]), .ip2(n22013), .op(n18769) );
  nand2_1 U21264 ( .ip1(n22014), .ip2(n18794), .op(n18768) );
  nand2_1 U21265 ( .ip1(n18769), .ip2(n18768), .op(n9904) );
  nand2_1 U21266 ( .ip1(\pipeline/csr/from_host [24]), .ip2(n22372), .op(
        n18771) );
  nand2_1 U21267 ( .ip1(n22373), .ip2(n18794), .op(n18770) );
  nand2_1 U21268 ( .ip1(n18771), .ip2(n18770), .op(n9936) );
  nand2_1 U21269 ( .ip1(n22378), .ip2(n18794), .op(n18773) );
  nand2_1 U21270 ( .ip1(\pipeline/csr/to_host [24]), .ip2(n22376), .op(n18772)
         );
  nand2_1 U21271 ( .ip1(n18773), .ip2(n18772), .op(n8748) );
  or2_1 U21272 ( .ip1(\pipeline/csr/cycle_full [24]), .ip2(n20136), .op(n18774) );
  nand2_1 U21273 ( .ip1(n18811), .ip2(n18774), .op(n18775) );
  or2_1 U21274 ( .ip1(n21145), .ip2(n18775), .op(n18777) );
  nand2_1 U21275 ( .ip1(n22021), .ip2(n18794), .op(n18776) );
  nand2_1 U21276 ( .ip1(n18777), .ip2(n18776), .op(\pipeline/csr/N1897 ) );
  nand2_1 U21277 ( .ip1(\pipeline/csr/mtimecmp [24]), .ip2(n22363), .op(n18779) );
  nand2_1 U21278 ( .ip1(n22365), .ip2(n18794), .op(n18778) );
  nand2_1 U21279 ( .ip1(n18779), .ip2(n18778), .op(n9998) );
  inv_1 U21280 ( .ip(n22274), .op(n22299) );
  nor2_1 U21281 ( .ip1(n22299), .ip2(n21001), .op(n18784) );
  inv_1 U21282 ( .ip(n18785), .op(n18782) );
  nor2_1 U21283 ( .ip1(\pipeline/csr/instret_full [23]), .ip2(n18780), .op(
        n18781) );
  nor3_1 U21284 ( .ip1(n21005), .ip2(n18782), .ip3(n18781), .op(n18783) );
  ab_or_c_or_d U21285 ( .ip1(n21016), .ip2(\pipeline/csr/instret_full [23]), 
        .ip3(n18784), .ip4(n18783), .op(n10115) );
  mux2_1 U21286 ( .ip1(\pipeline/csr/instret_full [24]), .ip2(n18786), .s(
        n18785), .op(n18787) );
  nor2_1 U21287 ( .ip1(n18787), .ip2(n18555), .op(n18789) );
  nor2_1 U21288 ( .ip1(n18787), .ip2(n21010), .op(n18788) );
  not_ab_or_c_or_d U21289 ( .ip1(n21016), .ip2(\pipeline/csr/instret_full [24]), .ip3(n18789), .ip4(n18788), .op(n18791) );
  nand2_1 U21290 ( .ip1(n21019), .ip2(n18794), .op(n18790) );
  nand2_1 U21291 ( .ip1(n18791), .ip2(n18790), .op(n10114) );
  nand2_1 U21292 ( .ip1(\pipeline/csr/mie [24]), .ip2(n22356), .op(n18793) );
  nand2_1 U21293 ( .ip1(n22357), .ip2(n18794), .op(n18792) );
  nand2_1 U21294 ( .ip1(n18793), .ip2(n18792), .op(n10036) );
  nand2_1 U21295 ( .ip1(n22314), .ip2(n18794), .op(n18797) );
  or2_1 U21296 ( .ip1(\pipeline/csr/cycle_full [56]), .ip2(n22300), .op(n18795) );
  nand3_1 U21297 ( .ip1(n18795), .ip2(n22309), .ip3(n22316), .op(n18796) );
  nand2_1 U21298 ( .ip1(n18797), .ip2(n18796), .op(\pipeline/csr/N1929 ) );
  nor2_1 U21299 ( .ip1(n22212), .ip2(n21110), .op(n18801) );
  inv_1 U21300 ( .ip(\pipeline/csr/instret_full [56]), .op(n18799) );
  nor2_1 U21301 ( .ip1(n18799), .ip2(n18798), .op(n18802) );
  not_ab_or_c_or_d U21302 ( .ip1(n18799), .ip2(n18798), .ip3(n18802), .ip4(
        n21111), .op(n18800) );
  ab_or_c_or_d U21303 ( .ip1(\pipeline/csr/instret_full [56]), .ip2(n21117), 
        .ip3(n18801), .ip4(n18800), .op(n10082) );
  nand2_1 U21304 ( .ip1(n20844), .ip2(n22217), .op(n18806) );
  nand2_1 U21305 ( .ip1(n21117), .ip2(\pipeline/csr/instret_full [57]), .op(
        n18805) );
  nand2_1 U21306 ( .ip1(\pipeline/csr/instret_full [57]), .ip2(n18802), .op(
        n19132) );
  or2_1 U21307 ( .ip1(\pipeline/csr/instret_full [57]), .ip2(n18802), .op(
        n18803) );
  nand3_1 U21308 ( .ip1(n20334), .ip2(n19132), .ip3(n18803), .op(n18804) );
  nand3_1 U21309 ( .ip1(n18806), .ip2(n18805), .ip3(n18804), .op(n10081) );
  nand2_1 U21310 ( .ip1(n22008), .ip2(n22217), .op(n18810) );
  xor2_1 U21311 ( .ip1(\pipeline/csr/mtime_full [25]), .ip2(n18807), .op(
        n18808) );
  nand2_1 U21312 ( .ip1(n18808), .ip2(n22009), .op(n18809) );
  nand2_1 U21313 ( .ip1(n18810), .ip2(n18809), .op(\pipeline/csr/N2106 ) );
  inv_1 U21314 ( .ip(n18811), .op(n18812) );
  nor2_1 U21315 ( .ip1(\pipeline/csr/cycle_full [25]), .ip2(n18812), .op(
        n18814) );
  nor3_1 U21316 ( .ip1(n19115), .ip2(n18814), .ip3(n21215), .op(n18813) );
  not_ab_or_c_or_d U21317 ( .ip1(n21076), .ip2(n22217), .ip3(n21217), .ip4(
        n18813), .op(n18817) );
  nor2_1 U21318 ( .ip1(n18814), .ip2(n19115), .op(n18815) );
  nor2_1 U21319 ( .ip1(n21198), .ip2(n18815), .op(n18816) );
  nor2_1 U21320 ( .ip1(n18817), .ip2(n18816), .op(\pipeline/csr/N1898 ) );
  inv_1 U21321 ( .ip(\pipeline/csr/instret_full [25]), .op(n18819) );
  nor2_1 U21322 ( .ip1(n18819), .ip2(n20990), .op(n18822) );
  mux2_1 U21323 ( .ip1(n18819), .ip2(\pipeline/csr/instret_full [25]), .s(
        n18818), .op(n18820) );
  nor2_1 U21324 ( .ip1(n21005), .ip2(n18820), .op(n18821) );
  ab_or_c_or_d U21325 ( .ip1(n21019), .ip2(n22217), .ip3(n18822), .ip4(n18821), 
        .op(n10113) );
  inv_1 U21326 ( .ip(n22217), .op(n22306) );
  nor2_1 U21327 ( .ip1(n22306), .ip2(n22267), .op(n18826) );
  not_ab_or_c_or_d U21328 ( .ip1(n18824), .ip2(n18823), .ip3(n19093), .ip4(
        n22276), .op(n18825) );
  or2_1 U21329 ( .ip1(n18826), .ip2(n18825), .op(\pipeline/csr/N1994 ) );
  nor2_1 U21330 ( .ip1(n22306), .ip2(n21168), .op(n18832) );
  inv_1 U21331 ( .ip(\pipeline/PC_WB [25]), .op(n18830) );
  inv_1 U21332 ( .ip(n18827), .op(n18828) );
  nand2_1 U21333 ( .ip1(n18828), .ip2(\pipeline/PC_WB [24]), .op(n18829) );
  not_ab_or_c_or_d U21334 ( .ip1(n18830), .ip2(n18829), .ip3(n19080), .ip4(
        n21171), .op(n18831) );
  ab_or_c_or_d U21335 ( .ip1(n21174), .ip2(\pipeline/epc [25]), .ip3(n18832), 
        .ip4(n18831), .op(n8846) );
  nand2_1 U21336 ( .ip1(n21995), .ip2(imem_haddr[27]), .op(n18834) );
  nand2_1 U21337 ( .ip1(\pipeline/PC_IF [27]), .ip2(n21996), .op(n18833) );
  nand2_1 U21338 ( .ip1(n18834), .ip2(n18833), .op(n8436) );
  nand2_1 U21339 ( .ip1(\pipeline/PC_IF [27]), .ip2(n22048), .op(n18836) );
  nand2_1 U21340 ( .ip1(\pipeline/PC_DX [27]), .ip2(n21999), .op(n18835) );
  nand2_1 U21341 ( .ip1(n18836), .ip2(n18835), .op(n8435) );
  nor2_1 U21342 ( .ip1(n18838), .ip2(n18837), .op(n21672) );
  nor2_1 U21343 ( .ip1(\pipeline/md_resp_result [27]), .ip2(n18839), .op(
        n18840) );
  nor2_1 U21344 ( .ip1(n18841), .ip2(n18840), .op(n18842) );
  nor2_1 U21345 ( .ip1(\pipeline/md/b [28]), .ip2(n18842), .op(n19026) );
  inv_1 U21346 ( .ip(n18842), .op(n18843) );
  nor2_1 U21347 ( .ip1(n18844), .ip2(n18843), .op(n19025) );
  nor2_1 U21348 ( .ip1(\pipeline/md_resp_result [28]), .ip2(n19025), .op(
        n18845) );
  nor2_1 U21349 ( .ip1(n19026), .ip2(n18845), .op(n18846) );
  nor2_1 U21350 ( .ip1(\pipeline/md/b [29]), .ip2(n18846), .op(n20682) );
  and2_1 U21351 ( .ip1(\pipeline/md/b [29]), .ip2(n18846), .op(n20681) );
  nor2_1 U21352 ( .ip1(\pipeline/md_resp_result [29]), .ip2(n20681), .op(
        n18847) );
  nor2_1 U21353 ( .ip1(n20682), .ip2(n18847), .op(n18848) );
  nor2_1 U21354 ( .ip1(\pipeline/md/b [30]), .ip2(n18848), .op(n21654) );
  inv_1 U21355 ( .ip(n18848), .op(n18849) );
  nor2_1 U21356 ( .ip1(n18850), .ip2(n18849), .op(n21652) );
  nor4_1 U21357 ( .ip1(\pipeline/md_resp_result [30]), .ip2(n21654), .ip3(
        n21652), .ip4(n22755), .op(n18861) );
  inv_1 U21358 ( .ip(n19017), .op(n19018) );
  nor2_1 U21359 ( .ip1(\pipeline/md/result [60]), .ip2(n19018), .op(n20672) );
  inv_1 U21360 ( .ip(\pipeline/md/result [61]), .op(n22743) );
  nand2_1 U21361 ( .ip1(n20672), .ip2(n22743), .op(n18851) );
  nor2_1 U21362 ( .ip1(\pipeline/md/result [62]), .ip2(n18851), .op(n21660) );
  not_ab_or_c_or_d U21363 ( .ip1(\pipeline/md/result [62]), .ip2(n18851), 
        .ip3(n21660), .ip4(n21505), .op(n18858) );
  inv_1 U21364 ( .ip(n18852), .op(n18853) );
  nor2_1 U21365 ( .ip1(n18853), .ip2(n21659), .op(n18856) );
  nor2_1 U21366 ( .ip1(n18856), .ip2(n18855), .op(n18854) );
  not_ab_or_c_or_d U21367 ( .ip1(n18856), .ip2(n18855), .ip3(n21960), .ip4(
        n18854), .op(n18857) );
  not_ab_or_c_or_d U21368 ( .ip1(\pipeline/md/result [62]), .ip2(n21509), 
        .ip3(n18858), .ip4(n18857), .op(n18859) );
  nor2_1 U21369 ( .ip1(n18859), .ip2(n21967), .op(n18860) );
  not_ab_or_c_or_d U21370 ( .ip1(n20306), .ip2(n21672), .ip3(n18861), .ip4(
        n18860), .op(n18866) );
  or2_1 U21371 ( .ip1(n21654), .ip2(n21652), .op(n18862) );
  nand2_1 U21372 ( .ip1(n20310), .ip2(n18862), .op(n18863) );
  nand2_1 U21373 ( .ip1(n22738), .ip2(n18863), .op(n18864) );
  nand2_1 U21374 ( .ip1(\pipeline/md_resp_result [30]), .ip2(n18864), .op(
        n18865) );
  nand2_1 U21375 ( .ip1(n18866), .ip2(n18865), .op(n8604) );
  mux2_1 U21376 ( .ip1(\pipeline/PC_WB [30]), .ip2(\pipeline/PC_DX [30]), .s(
        n17429), .op(n8873) );
  mux2_1 U21377 ( .ip1(\pipeline/PC_WB [27]), .ip2(\pipeline/PC_DX [27]), .s(
        n20389), .op(n8876) );
  mux2_1 U21378 ( .ip1(\pipeline/PC_WB [28]), .ip2(\pipeline/PC_DX [28]), .s(
        n22067), .op(n8875) );
  mux2_1 U21379 ( .ip1(\pipeline/PC_WB [26]), .ip2(\pipeline/PC_DX [26]), .s(
        n19498), .op(n8877) );
  nand2_1 U21380 ( .ip1(n18867), .ip2(n21583), .op(n18869) );
  nand2_1 U21381 ( .ip1(dmem_rdata[30]), .ip2(n21585), .op(n18868) );
  nand3_1 U21382 ( .ip1(n21588), .ip2(n18869), .ip3(n18868), .op(n18870) );
  mux2_1 U21383 ( .ip1(\pipeline/regfile/data[22][30] ), .ip2(n18870), .s(
        n19355), .op(n9194) );
  mux2_1 U21384 ( .ip1(\pipeline/regfile/data[28][30] ), .ip2(n18870), .s(
        n19359), .op(n9002) );
  mux2_1 U21385 ( .ip1(\pipeline/regfile/data[12][30] ), .ip2(n18870), .s(
        n19370), .op(n9514) );
  mux2_1 U21386 ( .ip1(\pipeline/regfile/data[19][30] ), .ip2(n18870), .s(
        n19361), .op(n9290) );
  mux2_1 U21387 ( .ip1(\pipeline/regfile/data[11][30] ), .ip2(n18870), .s(
        n19365), .op(n9546) );
  mux2_1 U21388 ( .ip1(\pipeline/regfile/data[30][30] ), .ip2(n18870), .s(
        n19363), .op(n8938) );
  mux2_1 U21389 ( .ip1(\pipeline/regfile/data[18][30] ), .ip2(n18870), .s(
        n19364), .op(n9322) );
  mux2_1 U21390 ( .ip1(\pipeline/regfile/data[23][30] ), .ip2(n18870), .s(
        n19369), .op(n9162) );
  mux2_1 U21391 ( .ip1(\pipeline/regfile/data[6][30] ), .ip2(n18870), .s(
        n19362), .op(n9706) );
  mux2_1 U21392 ( .ip1(\pipeline/regfile/data[5][30] ), .ip2(n18870), .s(
        n19356), .op(n9738) );
  mux2_1 U21393 ( .ip1(\pipeline/regfile/data[3][30] ), .ip2(n18870), .s(
        n19380), .op(n9802) );
  mux2_1 U21394 ( .ip1(\pipeline/regfile/data[13][30] ), .ip2(n18870), .s(
        n19367), .op(n9482) );
  mux2_1 U21395 ( .ip1(\pipeline/regfile/data[20][30] ), .ip2(n18870), .s(
        n19377), .op(n9258) );
  mux2_1 U21396 ( .ip1(\pipeline/regfile/data[25][30] ), .ip2(n18870), .s(
        n19366), .op(n9098) );
  mux2_1 U21397 ( .ip1(\pipeline/regfile/data[24][30] ), .ip2(n18870), .s(
        n19376), .op(n9130) );
  mux2_1 U21398 ( .ip1(\pipeline/regfile/data[14][30] ), .ip2(n18870), .s(
        n19354), .op(n9450) );
  mux2_1 U21399 ( .ip1(\pipeline/regfile/data[4][30] ), .ip2(n18870), .s(
        n19383), .op(n9770) );
  mux2_1 U21400 ( .ip1(\pipeline/regfile/data[31][30] ), .ip2(n18870), .s(
        n19360), .op(n8906) );
  mux2_1 U21401 ( .ip1(\pipeline/regfile/data[26][30] ), .ip2(n18870), .s(
        n19358), .op(n9066) );
  mux2_1 U21402 ( .ip1(\pipeline/regfile/data[16][30] ), .ip2(n18870), .s(
        n19379), .op(n9386) );
  mux2_1 U21403 ( .ip1(\pipeline/regfile/data[9][30] ), .ip2(n18870), .s(
        n19378), .op(n9610) );
  mux2_1 U21404 ( .ip1(\pipeline/regfile/data[2][30] ), .ip2(n18870), .s(
        n19382), .op(n9834) );
  mux2_1 U21405 ( .ip1(\pipeline/regfile/data[1][30] ), .ip2(n18870), .s(
        n19381), .op(n9866) );
  mux2_1 U21406 ( .ip1(\pipeline/regfile/data[27][30] ), .ip2(n18870), .s(
        n19357), .op(n9034) );
  mux2_1 U21407 ( .ip1(\pipeline/regfile/data[15][30] ), .ip2(n18870), .s(
        n19373), .op(n9418) );
  mux2_1 U21408 ( .ip1(\pipeline/regfile/data[7][30] ), .ip2(n18870), .s(
        n19371), .op(n9674) );
  mux2_1 U21409 ( .ip1(\pipeline/regfile/data[21][30] ), .ip2(n18870), .s(
        n19375), .op(n9226) );
  mux2_1 U21410 ( .ip1(\pipeline/regfile/data[17][30] ), .ip2(n18870), .s(
        n19368), .op(n9354) );
  mux2_1 U21411 ( .ip1(\pipeline/regfile/data[8][30] ), .ip2(n18870), .s(
        n19372), .op(n9642) );
  mux2_1 U21412 ( .ip1(\pipeline/regfile/data[10][30] ), .ip2(n18870), .s(
        n19374), .op(n9578) );
  mux2_1 U21413 ( .ip1(\pipeline/regfile/data[29][30] ), .ip2(n18870), .s(
        n19353), .op(n8970) );
  nor2_1 U21414 ( .ip1(n22258), .ip2(n21168), .op(n18875) );
  inv_1 U21415 ( .ip(\pipeline/PC_WB [30]), .op(n18873) );
  nand2_1 U21416 ( .ip1(n20320), .ip2(\pipeline/PC_WB [29]), .op(n18872) );
  nand3_1 U21417 ( .ip1(n20320), .ip2(\pipeline/PC_WB [29]), .ip3(
        \pipeline/PC_WB [30]), .op(n20847) );
  inv_1 U21418 ( .ip(n20847), .op(n18871) );
  not_ab_or_c_or_d U21419 ( .ip1(n18873), .ip2(n18872), .ip3(n18871), .ip4(
        n21171), .op(n18874) );
  ab_or_c_or_d U21420 ( .ip1(n21174), .ip2(\pipeline/epc [30]), .ip3(n18875), 
        .ip4(n18874), .op(n8841) );
  nor2_1 U21421 ( .ip1(n22313), .ip2(n21029), .op(n18879) );
  inv_1 U21422 ( .ip(\pipeline/csr/mtvec [30]), .op(n18876) );
  nor2_1 U21423 ( .ip1(n21089), .ip2(n18876), .op(n18877) );
  nor2_1 U21424 ( .ip1(n21032), .ip2(n18877), .op(n18878) );
  nor2_1 U21425 ( .ip1(n18879), .ip2(n18878), .op(n9962) );
  mux2_1 U21426 ( .ip1(dmem_haddr[30]), .ip2(\pipeline/alu_out_WB [30]), .s(
        n19505), .op(n8702) );
  nand2_1 U21427 ( .ip1(n22282), .ip2(n22313), .op(n18883) );
  or2_1 U21428 ( .ip1(\pipeline/csr/time_full [62]), .ip2(n18952), .op(n18880)
         );
  nand3_1 U21429 ( .ip1(n18881), .ip2(n18880), .ip3(n22284), .op(n18882) );
  nand2_1 U21430 ( .ip1(n18883), .ip2(n18882), .op(\pipeline/csr/N1999 ) );
  nor2_1 U21431 ( .ip1(n22234), .ip2(n21029), .op(n18887) );
  inv_1 U21432 ( .ip(\pipeline/csr/mtvec [29]), .op(n18884) );
  nor2_1 U21433 ( .ip1(n21089), .ip2(n18884), .op(n18885) );
  nor2_1 U21434 ( .ip1(n21032), .ip2(n18885), .op(n18886) );
  nor2_1 U21435 ( .ip1(n18887), .ip2(n18886), .op(n9963) );
  nand2_1 U21436 ( .ip1(\pipeline/csr/from_host [29]), .ip2(n22372), .op(
        n18889) );
  nand2_1 U21437 ( .ip1(n22373), .ip2(n22234), .op(n18888) );
  nand2_1 U21438 ( .ip1(n18889), .ip2(n18888), .op(n9931) );
  nand2_1 U21439 ( .ip1(n22378), .ip2(n22234), .op(n18891) );
  nand2_1 U21440 ( .ip1(\pipeline/csr/to_host [29]), .ip2(n22376), .op(n18890)
         );
  nand2_1 U21441 ( .ip1(n18891), .ip2(n18890), .op(n8743) );
  inv_1 U21442 ( .ip(n22234), .op(n18975) );
  nor2_1 U21443 ( .ip1(n18975), .ip2(n21001), .op(n18896) );
  nor2_1 U21444 ( .ip1(\pipeline/csr/instret_full [29]), .ip2(n18892), .op(
        n18893) );
  nor3_1 U21445 ( .ip1(n21005), .ip2(n18894), .ip3(n18893), .op(n18895) );
  ab_or_c_or_d U21446 ( .ip1(n21016), .ip2(\pipeline/csr/instret_full [29]), 
        .ip3(n18896), .ip4(n18895), .op(n10109) );
  nand2_1 U21447 ( .ip1(n22008), .ip2(n22234), .op(n18899) );
  xor2_1 U21448 ( .ip1(\pipeline/csr/mtime_full [29]), .ip2(n19265), .op(
        n18897) );
  nand2_1 U21449 ( .ip1(n18897), .ip2(n22009), .op(n18898) );
  nand2_1 U21450 ( .ip1(n18899), .ip2(n18898), .op(\pipeline/csr/N2110 ) );
  nand2_1 U21451 ( .ip1(\pipeline/csr/mscratch [29]), .ip2(n22013), .op(n18901) );
  nand2_1 U21452 ( .ip1(n22014), .ip2(n22234), .op(n18900) );
  nand2_1 U21453 ( .ip1(n18901), .ip2(n18900), .op(n9899) );
  nand2_1 U21454 ( .ip1(n18903), .ip2(n18902), .op(n18911) );
  inv_1 U21455 ( .ip(n19040), .op(n18906) );
  nor2_1 U21456 ( .ip1(n18904), .ip2(n17087), .op(n18905) );
  nor2_1 U21457 ( .ip1(n18906), .ip2(n18905), .op(n18909) );
  nand2_1 U21458 ( .ip1(n19042), .ip2(n19041), .op(n18907) );
  or2_1 U21459 ( .ip1(n18907), .ip2(n19177), .op(n18908) );
  nand2_1 U21460 ( .ip1(n18909), .ip2(n18908), .op(n18910) );
  xnor2_1 U21461 ( .ip1(n18911), .ip2(n18910), .op(n18912) );
  nand2_1 U21462 ( .ip1(n18912), .ip2(n21577), .op(n18951) );
  nand2_1 U21463 ( .ip1(n18914), .ip2(n18913), .op(n18915) );
  mux2_1 U21464 ( .ip1(n20905), .ip2(n18915), .s(n13881), .op(n18917) );
  nand2_1 U21465 ( .ip1(n18917), .ip2(n18916), .op(n20238) );
  nor2_1 U21466 ( .ip1(n19186), .ip2(n18918), .op(n20913) );
  nand2_1 U21467 ( .ip1(n20229), .ip2(n20913), .op(n18926) );
  nand2_1 U21468 ( .ip1(n10191), .ip2(n13600), .op(n18919) );
  nand2_1 U21469 ( .ip1(n18919), .ip2(n21557), .op(n18922) );
  nand3_1 U21470 ( .ip1(n20891), .ip2(n20904), .ip3(n18920), .op(n18921) );
  nand2_1 U21471 ( .ip1(n18922), .ip2(n18921), .op(n18923) );
  not_ab_or_c_or_d U21472 ( .ip1(n20911), .ip2(n18924), .ip3(n19066), .ip4(
        n18923), .op(n18925) );
  nand2_1 U21473 ( .ip1(n18926), .ip2(n18925), .op(n18943) );
  nand2_1 U21474 ( .ip1(n18927), .ip2(n20891), .op(n18928) );
  and2_1 U21475 ( .ip1(n18928), .ip2(n19427), .op(n18931) );
  nand4_1 U21476 ( .ip1(n18932), .ip2(n18931), .ip3(n18930), .ip4(n18929), 
        .op(n18933) );
  nand2_1 U21477 ( .ip1(n18933), .ip2(n20900), .op(n18941) );
  nor2_1 U21478 ( .ip1(n20885), .ip2(n18934), .op(n18940) );
  nor2_1 U21479 ( .ip1(n18936), .ip2(n18935), .op(n18939) );
  nor2_1 U21480 ( .ip1(n20887), .ip2(n18937), .op(n18938) );
  not_ab_or_c_or_d U21481 ( .ip1(n19205), .ip2(n20238), .ip3(n18943), .ip4(
        n18942), .op(n18950) );
  nor2_1 U21482 ( .ip1(n18918), .ip2(n18944), .op(n18947) );
  nor2_1 U21483 ( .ip1(n13166), .ip2(n18945), .op(n18946) );
  not_ab_or_c_or_d U21484 ( .ip1(n21540), .ip2(n18948), .ip3(n18947), .ip4(
        n18946), .op(n20240) );
  nand2_1 U21485 ( .ip1(n20240), .ip2(n19213), .op(n18949) );
  nand3_1 U21486 ( .ip1(n18951), .ip2(n18950), .ip3(n18949), .op(
        dmem_haddr[29]) );
  mux2_1 U21487 ( .ip1(dmem_haddr[29]), .ip2(\pipeline/alu_out_WB [29]), .s(
        n19505), .op(n8703) );
  nor2_1 U21488 ( .ip1(n18975), .ip2(n22267), .op(n18955) );
  not_ab_or_c_or_d U21489 ( .ip1(n22286), .ip2(n18953), .ip3(n18952), .ip4(
        n22276), .op(n18954) );
  or2_1 U21490 ( .ip1(n18955), .ip2(n18954), .op(\pipeline/csr/N1998 ) );
  inv_1 U21491 ( .ip(n19256), .op(n18956) );
  nor2_1 U21492 ( .ip1(\pipeline/csr/time_full [29]), .ip2(n18956), .op(n18958) );
  nor3_1 U21493 ( .ip1(n21177), .ip2(n22251), .ip3(n18958), .op(n18957) );
  not_ab_or_c_or_d U21494 ( .ip1(n21179), .ip2(n22234), .ip3(n21217), .ip4(
        n18957), .op(n18961) );
  nor2_1 U21495 ( .ip1(n18958), .ip2(n22251), .op(n18959) );
  nor2_1 U21496 ( .ip1(n21198), .ip2(n18959), .op(n18960) );
  nor2_1 U21497 ( .ip1(n18961), .ip2(n18960), .op(\pipeline/csr/N1966 ) );
  inv_1 U21498 ( .ip(n19278), .op(n18962) );
  nor2_1 U21499 ( .ip1(\pipeline/csr/cycle_full [29]), .ip2(n18962), .op(
        n18964) );
  nor3_1 U21500 ( .ip1(n18998), .ip2(n18964), .ip3(n21215), .op(n18963) );
  not_ab_or_c_or_d U21501 ( .ip1(n21076), .ip2(n22234), .ip3(n21217), .ip4(
        n18963), .op(n18967) );
  nor2_1 U21502 ( .ip1(n18964), .ip2(n18998), .op(n18965) );
  nor2_1 U21503 ( .ip1(n21198), .ip2(n18965), .op(n18966) );
  nor2_1 U21504 ( .ip1(n18967), .ip2(n18966), .op(\pipeline/csr/N1902 ) );
  nand2_1 U21505 ( .ip1(\pipeline/csr/mtimecmp [29]), .ip2(n22363), .op(n18969) );
  nand2_1 U21506 ( .ip1(n22365), .ip2(n22234), .op(n18968) );
  nand2_1 U21507 ( .ip1(n18969), .ip2(n18968), .op(n9993) );
  nand2_1 U21508 ( .ip1(\pipeline/csr/mie [29]), .ip2(n22356), .op(n18971) );
  nand2_1 U21509 ( .ip1(n22357), .ip2(n22234), .op(n18970) );
  nand2_1 U21510 ( .ip1(n18971), .ip2(n18970), .op(n10031) );
  nor2_1 U21511 ( .ip1(n18975), .ip2(n22305), .op(n18974) );
  not_ab_or_c_or_d U21512 ( .ip1(n19296), .ip2(n18972), .ip3(n22315), .ip4(
        n22308), .op(n18973) );
  or2_1 U21513 ( .ip1(n18974), .ip2(n18973), .op(\pipeline/csr/N1934 ) );
  nor2_1 U21514 ( .ip1(n18975), .ip2(n21110), .op(n18978) );
  inv_1 U21515 ( .ip(\pipeline/csr/instret_full [60]), .op(n19251) );
  inv_1 U21516 ( .ip(\pipeline/csr/instret_full [58]), .op(n19133) );
  nor2_1 U21517 ( .ip1(n19133), .ip2(n19132), .op(n19244) );
  nand2_1 U21518 ( .ip1(\pipeline/csr/instret_full [59]), .ip2(n19244), .op(
        n19250) );
  nor2_1 U21519 ( .ip1(n19251), .ip2(n19250), .op(n19249) );
  and2_1 U21520 ( .ip1(\pipeline/csr/instret_full [61]), .ip2(n19249), .op(
        n18980) );
  nor2_1 U21521 ( .ip1(\pipeline/csr/instret_full [61]), .ip2(n19249), .op(
        n18976) );
  nor3_1 U21522 ( .ip1(n21111), .ip2(n18980), .ip3(n18976), .op(n18977) );
  ab_or_c_or_d U21523 ( .ip1(\pipeline/csr/instret_full [61]), .ip2(n21117), 
        .ip3(n18978), .ip4(n18977), .op(n10077) );
  nand2_1 U21524 ( .ip1(\pipeline/csr/instret_full [62]), .ip2(n18980), .op(
        n20920) );
  nand2_1 U21525 ( .ip1(n20334), .ip2(n20920), .op(n18979) );
  nand2_1 U21526 ( .ip1(n19134), .ip2(n18979), .op(n20923) );
  inv_1 U21527 ( .ip(n20920), .op(n18982) );
  inv_1 U21528 ( .ip(n18980), .op(n18981) );
  nor3_1 U21529 ( .ip1(n21111), .ip2(n18982), .ip3(n18981), .op(n18984) );
  nor2_1 U21530 ( .ip1(n22258), .ip2(n21110), .op(n18983) );
  ab_or_c_or_d U21531 ( .ip1(\pipeline/csr/instret_full [62]), .ip2(n20923), 
        .ip3(n18984), .ip4(n18983), .op(n10076) );
  inv_1 U21532 ( .ip(n18985), .op(n18986) );
  nor2_1 U21533 ( .ip1(\pipeline/csr/mtime_full [30]), .ip2(n18986), .op(
        n18988) );
  nor3_1 U21534 ( .ip1(n21193), .ip2(n18988), .ip3(n20935), .op(n18987) );
  not_ab_or_c_or_d U21535 ( .ip1(n21195), .ip2(n22313), .ip3(n21217), .ip4(
        n18987), .op(n18991) );
  nor2_1 U21536 ( .ip1(n18988), .ip2(n20935), .op(n18989) );
  nor2_1 U21537 ( .ip1(n21198), .ip2(n18989), .op(n18990) );
  nor2_1 U21538 ( .ip1(n18991), .ip2(n18990), .op(\pipeline/csr/N2111 ) );
  nand2_1 U21539 ( .ip1(\pipeline/csr/mscratch [30]), .ip2(n22013), .op(n18993) );
  nand2_1 U21540 ( .ip1(n22014), .ip2(n22313), .op(n18992) );
  nand2_1 U21541 ( .ip1(n18993), .ip2(n18992), .op(n9898) );
  nand2_1 U21542 ( .ip1(\pipeline/csr/from_host [30]), .ip2(n22372), .op(
        n18995) );
  nand2_1 U21543 ( .ip1(n22373), .ip2(n22313), .op(n18994) );
  nand2_1 U21544 ( .ip1(n18995), .ip2(n18994), .op(n9930) );
  nand2_1 U21545 ( .ip1(n22378), .ip2(n22313), .op(n18997) );
  nand2_1 U21546 ( .ip1(\pipeline/csr/to_host [30]), .ip2(n22376), .op(n18996)
         );
  nand2_1 U21547 ( .ip1(n18997), .ip2(n18996), .op(n8742) );
  or2_1 U21548 ( .ip1(\pipeline/csr/cycle_full [30]), .ip2(n18998), .op(n18999) );
  nand2_1 U21549 ( .ip1(n20945), .ip2(n18999), .op(n19000) );
  or2_1 U21550 ( .ip1(n21145), .ip2(n19000), .op(n19002) );
  nand2_1 U21551 ( .ip1(n22021), .ip2(n22313), .op(n19001) );
  nand2_1 U21552 ( .ip1(n19002), .ip2(n19001), .op(\pipeline/csr/N1903 ) );
  nand2_1 U21553 ( .ip1(\pipeline/csr/mtimecmp [30]), .ip2(n22363), .op(n19004) );
  nand2_1 U21554 ( .ip1(n22365), .ip2(n22313), .op(n19003) );
  nand2_1 U21555 ( .ip1(n19004), .ip2(n19003), .op(n9992) );
  nor2_1 U21556 ( .ip1(n22258), .ip2(n21001), .op(n19008) );
  not_ab_or_c_or_d U21557 ( .ip1(n19006), .ip2(n19005), .ip3(n20954), .ip4(
        n21005), .op(n19007) );
  ab_or_c_or_d U21558 ( .ip1(n21016), .ip2(\pipeline/csr/instret_full [30]), 
        .ip3(n19008), .ip4(n19007), .op(n10108) );
  nand2_1 U21559 ( .ip1(\pipeline/csr/mie [30]), .ip2(n22356), .op(n19010) );
  nand2_1 U21560 ( .ip1(n22357), .ip2(n22313), .op(n19009) );
  nand2_1 U21561 ( .ip1(n19010), .ip2(n19009), .op(n10030) );
  inv_1 U21562 ( .ip(n19011), .op(n19012) );
  mux2_1 U21563 ( .ip1(\pipeline/csr_rdata_WB [30]), .ip2(n19012), .s(n17777), 
        .op(n8776) );
  nor4_1 U21564 ( .ip1(\pipeline/md_resp_result [28]), .ip2(n19026), .ip3(
        n19025), .ip4(n22755), .op(n19024) );
  nand2_1 U21565 ( .ip1(\pipeline/md/negate_output ), .ip2(n19013), .op(n19015) );
  nor2_1 U21566 ( .ip1(n19016), .ip2(n19015), .op(n19014) );
  not_ab_or_c_or_d U21567 ( .ip1(n19016), .ip2(n19015), .ip3(n21960), .ip4(
        n19014), .op(n19022) );
  nor3_1 U21568 ( .ip1(\pipeline/md/result [60]), .ip2(n21966), .ip3(n19017), 
        .op(n19020) );
  inv_1 U21569 ( .ip(\pipeline/md/result [60]), .op(n22733) );
  not_ab_or_c_or_d U21570 ( .ip1(\pipeline/md/negate_output ), .ip2(n19018), 
        .ip3(n21967), .ip4(n22733), .op(n19019) );
  nor3_1 U21571 ( .ip1(n21972), .ip2(n19020), .ip3(n19019), .op(n19021) );
  nor2_1 U21572 ( .ip1(n19022), .ip2(n19021), .op(n19023) );
  not_ab_or_c_or_d U21573 ( .ip1(n21672), .ip2(n21977), .ip3(n19024), .ip4(
        n19023), .op(n19031) );
  or2_1 U21574 ( .ip1(n19026), .ip2(n19025), .op(n19027) );
  nand2_1 U21575 ( .ip1(n21440), .ip2(n19027), .op(n19028) );
  nand2_1 U21576 ( .ip1(n22738), .ip2(n19028), .op(n19029) );
  nand2_1 U21577 ( .ip1(\pipeline/md_resp_result [28]), .ip2(n19029), .op(
        n19030) );
  nand2_1 U21578 ( .ip1(n19031), .ip2(n19030), .op(n8606) );
  nand2_1 U21579 ( .ip1(n19032), .ip2(n21583), .op(n19034) );
  nand2_1 U21580 ( .ip1(dmem_rdata[28]), .ip2(n21585), .op(n19033) );
  nand3_1 U21581 ( .ip1(n21588), .ip2(n19034), .ip3(n19033), .op(n19035) );
  mux2_1 U21582 ( .ip1(\pipeline/regfile/data[22][28] ), .ip2(n19035), .s(
        n19355), .op(n9196) );
  mux2_1 U21583 ( .ip1(\pipeline/regfile/data[28][28] ), .ip2(n19035), .s(
        n19359), .op(n9004) );
  mux2_1 U21584 ( .ip1(\pipeline/regfile/data[12][28] ), .ip2(n19035), .s(
        n19370), .op(n9516) );
  mux2_1 U21585 ( .ip1(\pipeline/regfile/data[19][28] ), .ip2(n19035), .s(
        n19361), .op(n9292) );
  mux2_1 U21586 ( .ip1(\pipeline/regfile/data[11][28] ), .ip2(n19035), .s(
        n19365), .op(n9548) );
  mux2_1 U21587 ( .ip1(\pipeline/regfile/data[30][28] ), .ip2(n19035), .s(
        n19363), .op(n8940) );
  mux2_1 U21588 ( .ip1(\pipeline/regfile/data[18][28] ), .ip2(n19035), .s(
        n19364), .op(n9324) );
  mux2_1 U21589 ( .ip1(\pipeline/regfile/data[23][28] ), .ip2(n19035), .s(
        n19369), .op(n9164) );
  mux2_1 U21590 ( .ip1(\pipeline/regfile/data[6][28] ), .ip2(n19035), .s(
        n19362), .op(n9708) );
  mux2_1 U21591 ( .ip1(\pipeline/regfile/data[5][28] ), .ip2(n19035), .s(
        n19356), .op(n9740) );
  mux2_1 U21592 ( .ip1(\pipeline/regfile/data[3][28] ), .ip2(n19035), .s(
        n19380), .op(n9804) );
  mux2_1 U21593 ( .ip1(\pipeline/regfile/data[13][28] ), .ip2(n19035), .s(
        n19367), .op(n9484) );
  mux2_1 U21594 ( .ip1(\pipeline/regfile/data[20][28] ), .ip2(n19035), .s(
        n19377), .op(n9260) );
  mux2_1 U21595 ( .ip1(\pipeline/regfile/data[25][28] ), .ip2(n19035), .s(
        n19366), .op(n9100) );
  mux2_1 U21596 ( .ip1(\pipeline/regfile/data[24][28] ), .ip2(n19035), .s(
        n19376), .op(n9132) );
  mux2_1 U21597 ( .ip1(\pipeline/regfile/data[14][28] ), .ip2(n19035), .s(
        n19354), .op(n9452) );
  mux2_1 U21598 ( .ip1(\pipeline/regfile/data[4][28] ), .ip2(n19035), .s(
        n19383), .op(n9772) );
  mux2_1 U21599 ( .ip1(\pipeline/regfile/data[31][28] ), .ip2(n19035), .s(
        n19360), .op(n8908) );
  mux2_1 U21600 ( .ip1(\pipeline/regfile/data[26][28] ), .ip2(n19035), .s(
        n19358), .op(n9068) );
  mux2_1 U21601 ( .ip1(\pipeline/regfile/data[16][28] ), .ip2(n19035), .s(
        n19379), .op(n9388) );
  mux2_1 U21602 ( .ip1(\pipeline/regfile/data[9][28] ), .ip2(n19035), .s(
        n19378), .op(n9612) );
  mux2_1 U21603 ( .ip1(\pipeline/regfile/data[2][28] ), .ip2(n19035), .s(
        n19382), .op(n9836) );
  mux2_1 U21604 ( .ip1(\pipeline/regfile/data[1][28] ), .ip2(n19035), .s(
        n19381), .op(n9868) );
  mux2_1 U21605 ( .ip1(\pipeline/regfile/data[27][28] ), .ip2(n19035), .s(
        n19357), .op(n9036) );
  mux2_1 U21606 ( .ip1(\pipeline/regfile/data[15][28] ), .ip2(n19035), .s(
        n19373), .op(n9420) );
  mux2_1 U21607 ( .ip1(\pipeline/regfile/data[7][28] ), .ip2(n19035), .s(
        n19371), .op(n9676) );
  mux2_1 U21608 ( .ip1(\pipeline/regfile/data[21][28] ), .ip2(n19035), .s(
        n19375), .op(n9228) );
  mux2_1 U21609 ( .ip1(\pipeline/regfile/data[17][28] ), .ip2(n19035), .s(
        n19368), .op(n9356) );
  mux2_1 U21610 ( .ip1(\pipeline/regfile/data[8][28] ), .ip2(n19035), .s(
        n19372), .op(n9644) );
  mux2_1 U21611 ( .ip1(\pipeline/regfile/data[10][28] ), .ip2(n19035), .s(
        n19374), .op(n9580) );
  mux2_1 U21612 ( .ip1(\pipeline/regfile/data[29][28] ), .ip2(n19035), .s(
        n19353), .op(n8972) );
  nor2_1 U21613 ( .ip1(n22281), .ip2(n21029), .op(n19039) );
  inv_1 U21614 ( .ip(\pipeline/csr/mtvec [28]), .op(n19036) );
  nor2_1 U21615 ( .ip1(n21089), .ip2(n19036), .op(n19037) );
  nor2_1 U21616 ( .ip1(n21032), .ip2(n19037), .op(n19038) );
  nor2_1 U21617 ( .ip1(n19039), .ip2(n19038), .op(n9964) );
  nand2_1 U21618 ( .ip1(n19041), .ip2(n19040), .op(n19045) );
  nand2_1 U21619 ( .ip1(n20878), .ip2(n19042), .op(n19043) );
  nand2_1 U21620 ( .ip1(n17087), .ip2(n19043), .op(n19044) );
  xnor2_1 U21621 ( .ip1(n19045), .ip2(n19044), .op(n19079) );
  nor2_1 U21622 ( .ip1(n18918), .ip2(n19046), .op(n19049) );
  nor2_1 U21623 ( .ip1(n13881), .ip2(n19047), .op(n19048) );
  ab_or_c_or_d U21624 ( .ip1(n21540), .ip2(n19050), .ip3(n19049), .ip4(n19048), 
        .op(n20723) );
  nor2_1 U21625 ( .ip1(n20883), .ip2(n20723), .op(n19078) );
  nor2_1 U21626 ( .ip1(n10180), .ip2(n21532), .op(n19055) );
  nand2_1 U21627 ( .ip1(n20892), .ip2(n19199), .op(n19053) );
  nand2_1 U21628 ( .ip1(n21536), .ip2(n19051), .op(n19052) );
  nand3_1 U21629 ( .ip1(n19053), .ip2(n19052), .ip3(n19427), .op(n19054) );
  not_ab_or_c_or_d U21630 ( .ip1(n19056), .ip2(n13651), .ip3(n19055), .ip4(
        n19054), .op(n19057) );
  not_ab_or_c_or_d U21631 ( .ip1(n21540), .ip2(n19058), .ip3(n19057), .ip4(
        n20724), .op(n19063) );
  nand2_1 U21632 ( .ip1(n19059), .ip2(n20896), .op(n19062) );
  nand2_1 U21633 ( .ip1(n19060), .ip2(n19193), .op(n19061) );
  nand3_1 U21634 ( .ip1(n19063), .ip2(n19062), .ip3(n19061), .op(n19076) );
  nor2_1 U21635 ( .ip1(n19427), .ip2(n19064), .op(n19065) );
  nor2_1 U21636 ( .ip1(n19066), .ip2(n19065), .op(n19208) );
  nor3_1 U21637 ( .ip1(n19067), .ip2(n21551), .ip3(n10180), .op(n19072) );
  nor2_1 U21638 ( .ip1(n19069), .ip2(n19068), .op(n19070) );
  nor2_1 U21639 ( .ip1(n20907), .ip2(n19070), .op(n19071) );
  not_ab_or_c_or_d U21640 ( .ip1(n20911), .ip2(n19073), .ip3(n19072), .ip4(
        n19071), .op(n19075) );
  nand3_1 U21641 ( .ip1(n20733), .ip2(n19427), .ip3(n21572), .op(n19074) );
  nand4_1 U21642 ( .ip1(n19076), .ip2(n19208), .ip3(n19075), .ip4(n19074), 
        .op(n19077) );
  ab_or_c_or_d U21643 ( .ip1(n19079), .ip2(n21577), .ip3(n19078), .ip4(n19077), 
        .op(dmem_haddr[28]) );
  mux2_1 U21644 ( .ip1(dmem_haddr[28]), .ip2(\pipeline/alu_out_WB [28]), .s(
        n19505), .op(n8704) );
  nand2_1 U21645 ( .ip1(n21043), .ip2(n22222), .op(n19084) );
  xor2_1 U21646 ( .ip1(n19080), .ip2(\pipeline/PC_WB [26]), .op(n19081) );
  nand2_1 U21647 ( .ip1(n21046), .ip2(n19081), .op(n19083) );
  nand2_1 U21648 ( .ip1(\pipeline/epc [26]), .ip2(n21174), .op(n19082) );
  nand3_1 U21649 ( .ip1(n19084), .ip2(n19083), .ip3(n19082), .op(n8845) );
  nor2_1 U21650 ( .ip1(n22222), .ip2(n21029), .op(n19088) );
  inv_1 U21651 ( .ip(\pipeline/csr/mtvec [26]), .op(n19085) );
  nor2_1 U21652 ( .ip1(n21089), .ip2(n19085), .op(n19086) );
  nor2_1 U21653 ( .ip1(n21032), .ip2(n19086), .op(n19087) );
  nor2_1 U21654 ( .ip1(n19088), .ip2(n19087), .op(n9966) );
  nand2_1 U21655 ( .ip1(n19089), .ip2(n21583), .op(n19091) );
  nand2_1 U21656 ( .ip1(n21585), .ip2(dmem_rdata[26]), .op(n19090) );
  nand3_1 U21657 ( .ip1(n21588), .ip2(n19091), .ip3(n19090), .op(n19092) );
  mux2_1 U21658 ( .ip1(\pipeline/regfile/data[29][26] ), .ip2(n19092), .s(
        n19353), .op(n8974) );
  mux2_1 U21659 ( .ip1(\pipeline/regfile/data[14][26] ), .ip2(n19092), .s(
        n19354), .op(n9454) );
  mux2_1 U21660 ( .ip1(\pipeline/regfile/data[22][26] ), .ip2(n19092), .s(
        n19355), .op(n9198) );
  mux2_1 U21661 ( .ip1(\pipeline/regfile/data[5][26] ), .ip2(n19092), .s(
        n19356), .op(n9742) );
  mux2_1 U21662 ( .ip1(\pipeline/regfile/data[27][26] ), .ip2(n19092), .s(
        n19357), .op(n9038) );
  mux2_1 U21663 ( .ip1(\pipeline/regfile/data[26][26] ), .ip2(n19092), .s(
        n19358), .op(n9070) );
  mux2_1 U21664 ( .ip1(\pipeline/regfile/data[28][26] ), .ip2(n19092), .s(
        n19359), .op(n9006) );
  mux2_1 U21665 ( .ip1(\pipeline/regfile/data[31][26] ), .ip2(n19092), .s(
        n19360), .op(n8910) );
  mux2_1 U21666 ( .ip1(\pipeline/regfile/data[19][26] ), .ip2(n19092), .s(
        n19361), .op(n9294) );
  mux2_1 U21667 ( .ip1(\pipeline/regfile/data[6][26] ), .ip2(n19092), .s(
        n19362), .op(n9710) );
  mux2_1 U21668 ( .ip1(\pipeline/regfile/data[30][26] ), .ip2(n19092), .s(
        n19363), .op(n8942) );
  mux2_1 U21669 ( .ip1(\pipeline/regfile/data[18][26] ), .ip2(n19092), .s(
        n19364), .op(n9326) );
  mux2_1 U21670 ( .ip1(\pipeline/regfile/data[11][26] ), .ip2(n19092), .s(
        n19365), .op(n9550) );
  mux2_1 U21671 ( .ip1(\pipeline/regfile/data[25][26] ), .ip2(n19092), .s(
        n19366), .op(n9102) );
  mux2_1 U21672 ( .ip1(\pipeline/regfile/data[13][26] ), .ip2(n19092), .s(
        n19367), .op(n9486) );
  mux2_1 U21673 ( .ip1(\pipeline/regfile/data[17][26] ), .ip2(n19092), .s(
        n19368), .op(n9358) );
  mux2_1 U21674 ( .ip1(\pipeline/regfile/data[23][26] ), .ip2(n19092), .s(
        n19369), .op(n9166) );
  mux2_1 U21675 ( .ip1(\pipeline/regfile/data[12][26] ), .ip2(n19092), .s(
        n19370), .op(n9518) );
  mux2_1 U21676 ( .ip1(\pipeline/regfile/data[7][26] ), .ip2(n19092), .s(
        n19371), .op(n9678) );
  mux2_1 U21677 ( .ip1(\pipeline/regfile/data[8][26] ), .ip2(n19092), .s(
        n19372), .op(n9646) );
  mux2_1 U21678 ( .ip1(\pipeline/regfile/data[15][26] ), .ip2(n19092), .s(
        n19373), .op(n9422) );
  mux2_1 U21679 ( .ip1(\pipeline/regfile/data[10][26] ), .ip2(n19092), .s(
        n19374), .op(n9582) );
  mux2_1 U21680 ( .ip1(\pipeline/regfile/data[21][26] ), .ip2(n19092), .s(
        n19375), .op(n9230) );
  mux2_1 U21681 ( .ip1(\pipeline/regfile/data[24][26] ), .ip2(n19092), .s(
        n19376), .op(n9134) );
  mux2_1 U21682 ( .ip1(\pipeline/regfile/data[20][26] ), .ip2(n19092), .s(
        n19377), .op(n9262) );
  mux2_1 U21683 ( .ip1(\pipeline/regfile/data[9][26] ), .ip2(n19092), .s(
        n19378), .op(n9614) );
  mux2_1 U21684 ( .ip1(\pipeline/regfile/data[16][26] ), .ip2(n19092), .s(
        n19379), .op(n9390) );
  mux2_1 U21685 ( .ip1(\pipeline/regfile/data[3][26] ), .ip2(n19092), .s(
        n19380), .op(n9806) );
  mux2_1 U21686 ( .ip1(\pipeline/regfile/data[1][26] ), .ip2(n19092), .s(
        n19381), .op(n9870) );
  mux2_1 U21687 ( .ip1(\pipeline/regfile/data[2][26] ), .ip2(n19092), .s(
        n19382), .op(n9838) );
  mux2_1 U21688 ( .ip1(\pipeline/regfile/data[4][26] ), .ip2(n19092), .s(
        n19383), .op(n9774) );
  mux2_1 U21689 ( .ip1(dmem_haddr[26]), .ip2(\pipeline/alu_out_WB [26]), .s(
        n19505), .op(n8706) );
  nand2_1 U21690 ( .ip1(n22282), .ip2(n22222), .op(n19096) );
  or2_1 U21691 ( .ip1(\pipeline/csr/time_full [58]), .ip2(n19093), .op(n19094)
         );
  nand3_1 U21692 ( .ip1(n19239), .ip2(n19094), .ip3(n22284), .op(n19095) );
  nand2_1 U21693 ( .ip1(n19096), .ip2(n19095), .op(\pipeline/csr/N1995 ) );
  or2_1 U21694 ( .ip1(\pipeline/csr/time_full [26]), .ip2(n19097), .op(n19098)
         );
  nand2_1 U21695 ( .ip1(n19216), .ip2(n19098), .op(n19099) );
  or2_1 U21696 ( .ip1(n22002), .ip2(n19099), .op(n19101) );
  nand2_1 U21697 ( .ip1(n22005), .ip2(n22222), .op(n19100) );
  nand2_1 U21698 ( .ip1(n19101), .ip2(n19100), .op(\pipeline/csr/N1963 ) );
  inv_1 U21699 ( .ip(n19102), .op(n19103) );
  nor2_1 U21700 ( .ip1(\pipeline/csr/mtime_full [26]), .ip2(n19103), .op(
        n19105) );
  nor3_1 U21701 ( .ip1(n21193), .ip2(n19105), .ip3(n19155), .op(n19104) );
  not_ab_or_c_or_d U21702 ( .ip1(n21195), .ip2(n22222), .ip3(n21217), .ip4(
        n19104), .op(n19108) );
  nor2_1 U21703 ( .ip1(n19105), .ip2(n19155), .op(n19106) );
  nor2_1 U21704 ( .ip1(n21198), .ip2(n19106), .op(n19107) );
  nor2_1 U21705 ( .ip1(n19108), .ip2(n19107), .op(\pipeline/csr/N2107 ) );
  nand2_1 U21706 ( .ip1(\pipeline/csr/mscratch [26]), .ip2(n22013), .op(n19110) );
  nand2_1 U21707 ( .ip1(n22014), .ip2(n22222), .op(n19109) );
  nand2_1 U21708 ( .ip1(n19110), .ip2(n19109), .op(n9902) );
  nand2_1 U21709 ( .ip1(\pipeline/csr/from_host [26]), .ip2(n22372), .op(
        n19112) );
  nand2_1 U21710 ( .ip1(n22373), .ip2(n22222), .op(n19111) );
  nand2_1 U21711 ( .ip1(n19112), .ip2(n19111), .op(n9934) );
  nand2_1 U21712 ( .ip1(n22378), .ip2(n22222), .op(n19114) );
  nand2_1 U21713 ( .ip1(\pipeline/csr/to_host [26]), .ip2(n22376), .op(n19113)
         );
  nand2_1 U21714 ( .ip1(n19114), .ip2(n19113), .op(n8746) );
  or2_1 U21715 ( .ip1(\pipeline/csr/cycle_full [26]), .ip2(n19115), .op(n19116) );
  nand2_1 U21716 ( .ip1(n19223), .ip2(n19116), .op(n19117) );
  or2_1 U21717 ( .ip1(n21145), .ip2(n19117), .op(n19119) );
  nand2_1 U21718 ( .ip1(n22021), .ip2(n22222), .op(n19118) );
  nand2_1 U21719 ( .ip1(n19119), .ip2(n19118), .op(\pipeline/csr/N1899 ) );
  nand2_1 U21720 ( .ip1(\pipeline/csr/mtimecmp [26]), .ip2(n22363), .op(n19121) );
  nand2_1 U21721 ( .ip1(n22365), .ip2(n22222), .op(n19120) );
  nand2_1 U21722 ( .ip1(n19121), .ip2(n19120), .op(n9996) );
  mux2_1 U21723 ( .ip1(\pipeline/csr/instret_full [26]), .ip2(n19125), .s(
        n19122), .op(n19124) );
  nor2_1 U21724 ( .ip1(n21012), .ip2(n21011), .op(n19123) );
  nor2_1 U21725 ( .ip1(n19124), .ip2(n19123), .op(n19127) );
  nor2_1 U21726 ( .ip1(n19125), .ip2(n20990), .op(n19126) );
  nor2_1 U21727 ( .ip1(n19127), .ip2(n19126), .op(n19129) );
  nand2_1 U21728 ( .ip1(n21019), .ip2(n22222), .op(n19128) );
  nand2_1 U21729 ( .ip1(n19129), .ip2(n19128), .op(n10112) );
  nand2_1 U21730 ( .ip1(\pipeline/csr/mie [26]), .ip2(n22356), .op(n19131) );
  nand2_1 U21731 ( .ip1(n22357), .ip2(n22222), .op(n19130) );
  nand2_1 U21732 ( .ip1(n19131), .ip2(n19130), .op(n10034) );
  not_ab_or_c_or_d U21733 ( .ip1(n19133), .ip2(n19132), .ip3(n19244), .ip4(
        n21111), .op(n19136) );
  nor2_1 U21734 ( .ip1(n19134), .ip2(n19133), .op(n19135) );
  ab_or_c_or_d U21735 ( .ip1(n20844), .ip2(n22222), .ip3(n19136), .ip4(n19135), 
        .op(n10080) );
  nor2_1 U21736 ( .ip1(n19243), .ip2(n21029), .op(n19140) );
  inv_1 U21737 ( .ip(\pipeline/csr/mtvec [27]), .op(n19137) );
  nor2_1 U21738 ( .ip1(htif_reset), .ip2(n19137), .op(n19138) );
  nor2_1 U21739 ( .ip1(n21032), .ip2(n19138), .op(n19139) );
  nor2_1 U21740 ( .ip1(n19140), .ip2(n19139), .op(n9965) );
  nand2_1 U21741 ( .ip1(\pipeline/csr/from_host [27]), .ip2(n22372), .op(
        n19142) );
  nand2_1 U21742 ( .ip1(n22373), .ip2(n19243), .op(n19141) );
  nand2_1 U21743 ( .ip1(n19142), .ip2(n19141), .op(n9933) );
  nand2_1 U21744 ( .ip1(n22378), .ip2(n19243), .op(n19144) );
  nand2_1 U21745 ( .ip1(\pipeline/csr/to_host [27]), .ip2(n22376), .op(n19143)
         );
  nand2_1 U21746 ( .ip1(n19144), .ip2(n19143), .op(n8745) );
  inv_1 U21747 ( .ip(\pipeline/csr/instret_full [27]), .op(n19146) );
  nor2_1 U21748 ( .ip1(n19146), .ip2(n20990), .op(n19149) );
  mux2_1 U21749 ( .ip1(n19146), .ip2(\pipeline/csr/instret_full [27]), .s(
        n19145), .op(n19147) );
  nor2_1 U21750 ( .ip1(n21005), .ip2(n19147), .op(n19148) );
  ab_or_c_or_d U21751 ( .ip1(n21019), .ip2(n19243), .ip3(n19149), .ip4(n19148), 
        .op(n10111) );
  nand2_1 U21752 ( .ip1(n21043), .ip2(n19243), .op(n19154) );
  xor2_1 U21753 ( .ip1(n19150), .ip2(\pipeline/PC_WB [27]), .op(n19151) );
  nand2_1 U21754 ( .ip1(n21046), .ip2(n19151), .op(n19153) );
  nand2_1 U21755 ( .ip1(\pipeline/epc [27]), .ip2(n21174), .op(n19152) );
  nand3_1 U21756 ( .ip1(n19154), .ip2(n19153), .ip3(n19152), .op(n8844) );
  inv_1 U21757 ( .ip(\pipeline/csr/mtime_full [27]), .op(n19613) );
  xor2_1 U21758 ( .ip1(n19155), .ip2(n19613), .op(n19157) );
  nor2_1 U21759 ( .ip1(n21193), .ip2(n19157), .op(n19156) );
  not_ab_or_c_or_d U21760 ( .ip1(n21195), .ip2(n19243), .ip3(n21217), .ip4(
        n19156), .op(n19160) );
  inv_1 U21761 ( .ip(n19157), .op(n19158) );
  nor2_1 U21762 ( .ip1(n22254), .ip2(n19158), .op(n19159) );
  nor2_1 U21763 ( .ip1(n19160), .ip2(n19159), .op(\pipeline/csr/N2108 ) );
  nand2_1 U21764 ( .ip1(\pipeline/csr/mscratch [27]), .ip2(n22013), .op(n19162) );
  nand2_1 U21765 ( .ip1(n22014), .ip2(n19243), .op(n19161) );
  nand2_1 U21766 ( .ip1(n19162), .ip2(n19161), .op(n9901) );
  inv_1 U21767 ( .ip(n22244), .op(n22235) );
  nand2_1 U21768 ( .ip1(n22235), .ip2(n19243), .op(n19165) );
  inv_1 U21769 ( .ip(\pipeline/csr/mtime_full [56]), .op(n22214) );
  inv_1 U21770 ( .ip(\pipeline/csr/mtime_full [54]), .op(n22205) );
  nand2_1 U21771 ( .ip1(\pipeline/csr/mtime_full [51]), .ip2(n22190), .op(
        n22195) );
  nor2_1 U21772 ( .ip1(n22196), .ip2(n22195), .op(n22199) );
  nand2_1 U21773 ( .ip1(\pipeline/csr/mtime_full [53]), .ip2(n22199), .op(
        n22204) );
  nor2_1 U21774 ( .ip1(n22205), .ip2(n22204), .op(n22208) );
  nand2_1 U21775 ( .ip1(\pipeline/csr/mtime_full [55]), .ip2(n22208), .op(
        n22213) );
  nor2_1 U21776 ( .ip1(n22214), .ip2(n22213), .op(n22218) );
  nand2_1 U21777 ( .ip1(\pipeline/csr/mtime_full [57]), .ip2(n22218), .op(
        n22225) );
  nor2_1 U21778 ( .ip1(n22226), .ip2(n22225), .op(n22224) );
  or2_1 U21779 ( .ip1(\pipeline/csr/mtime_full [59]), .ip2(n22224), .op(n19163) );
  nand2_1 U21780 ( .ip1(\pipeline/csr/mtime_full [59]), .ip2(n22224), .op(
        n22230) );
  nand3_1 U21781 ( .ip1(n19163), .ip2(n22230), .ip3(n18449), .op(n19164) );
  nand2_1 U21782 ( .ip1(n19165), .ip2(n19164), .op(\pipeline/csr/N2140 ) );
  nand2_1 U21783 ( .ip1(n19166), .ip2(n21583), .op(n19168) );
  nand2_1 U21784 ( .ip1(dmem_rdata[27]), .ip2(n21585), .op(n19167) );
  nand3_1 U21785 ( .ip1(n21588), .ip2(n19168), .ip3(n19167), .op(n19169) );
  mux2_1 U21786 ( .ip1(\pipeline/regfile/data[29][27] ), .ip2(n19169), .s(
        n19353), .op(n8973) );
  mux2_1 U21787 ( .ip1(\pipeline/regfile/data[14][27] ), .ip2(n19169), .s(
        n19354), .op(n9453) );
  mux2_1 U21788 ( .ip1(\pipeline/regfile/data[22][27] ), .ip2(n19169), .s(
        n19355), .op(n9197) );
  mux2_1 U21789 ( .ip1(\pipeline/regfile/data[5][27] ), .ip2(n19169), .s(
        n19356), .op(n9741) );
  mux2_1 U21790 ( .ip1(\pipeline/regfile/data[27][27] ), .ip2(n19169), .s(
        n19357), .op(n9037) );
  mux2_1 U21791 ( .ip1(\pipeline/regfile/data[26][27] ), .ip2(n19169), .s(
        n19358), .op(n9069) );
  mux2_1 U21792 ( .ip1(\pipeline/regfile/data[28][27] ), .ip2(n19169), .s(
        n19359), .op(n9005) );
  mux2_1 U21793 ( .ip1(\pipeline/regfile/data[31][27] ), .ip2(n19169), .s(
        n19360), .op(n8909) );
  mux2_1 U21794 ( .ip1(\pipeline/regfile/data[19][27] ), .ip2(n19169), .s(
        n19361), .op(n9293) );
  mux2_1 U21795 ( .ip1(\pipeline/regfile/data[6][27] ), .ip2(n19169), .s(
        n19362), .op(n9709) );
  mux2_1 U21796 ( .ip1(\pipeline/regfile/data[30][27] ), .ip2(n19169), .s(
        n19363), .op(n8941) );
  mux2_1 U21797 ( .ip1(\pipeline/regfile/data[18][27] ), .ip2(n19169), .s(
        n19364), .op(n9325) );
  mux2_1 U21798 ( .ip1(\pipeline/regfile/data[11][27] ), .ip2(n19169), .s(
        n19365), .op(n9549) );
  mux2_1 U21799 ( .ip1(\pipeline/regfile/data[25][27] ), .ip2(n19169), .s(
        n19366), .op(n9101) );
  mux2_1 U21800 ( .ip1(\pipeline/regfile/data[13][27] ), .ip2(n19169), .s(
        n19367), .op(n9485) );
  mux2_1 U21801 ( .ip1(\pipeline/regfile/data[17][27] ), .ip2(n19169), .s(
        n19368), .op(n9357) );
  mux2_1 U21802 ( .ip1(\pipeline/regfile/data[23][27] ), .ip2(n19169), .s(
        n19369), .op(n9165) );
  mux2_1 U21803 ( .ip1(\pipeline/regfile/data[12][27] ), .ip2(n19169), .s(
        n19370), .op(n9517) );
  mux2_1 U21804 ( .ip1(\pipeline/regfile/data[7][27] ), .ip2(n19169), .s(
        n19371), .op(n9677) );
  mux2_1 U21805 ( .ip1(\pipeline/regfile/data[8][27] ), .ip2(n19169), .s(
        n19372), .op(n9645) );
  mux2_1 U21806 ( .ip1(\pipeline/regfile/data[15][27] ), .ip2(n19169), .s(
        n19373), .op(n9421) );
  mux2_1 U21807 ( .ip1(\pipeline/regfile/data[10][27] ), .ip2(n19169), .s(
        n19374), .op(n9581) );
  mux2_1 U21808 ( .ip1(\pipeline/regfile/data[21][27] ), .ip2(n19169), .s(
        n19375), .op(n9229) );
  mux2_1 U21809 ( .ip1(\pipeline/regfile/data[24][27] ), .ip2(n19169), .s(
        n19376), .op(n9133) );
  mux2_1 U21810 ( .ip1(\pipeline/regfile/data[20][27] ), .ip2(n19169), .s(
        n19377), .op(n9261) );
  mux2_1 U21811 ( .ip1(\pipeline/regfile/data[9][27] ), .ip2(n19169), .s(
        n19378), .op(n9613) );
  mux2_1 U21812 ( .ip1(\pipeline/regfile/data[16][27] ), .ip2(n19169), .s(
        n19379), .op(n9389) );
  mux2_1 U21813 ( .ip1(\pipeline/regfile/data[3][27] ), .ip2(n19169), .s(
        n19380), .op(n9805) );
  mux2_1 U21814 ( .ip1(\pipeline/regfile/data[1][27] ), .ip2(n19169), .s(
        n19381), .op(n9869) );
  mux2_1 U21815 ( .ip1(\pipeline/regfile/data[2][27] ), .ip2(n19169), .s(
        n19382), .op(n9837) );
  mux2_1 U21816 ( .ip1(\pipeline/regfile/data[4][27] ), .ip2(n19169), .s(
        n19383), .op(n9773) );
  nand2_1 U21817 ( .ip1(n19171), .ip2(n19170), .op(n19182) );
  nor2_1 U21818 ( .ip1(n20871), .ip2(n19172), .op(n19173) );
  nor2_1 U21819 ( .ip1(n19174), .ip2(n19173), .op(n19180) );
  nand2_1 U21820 ( .ip1(n19176), .ip2(n19175), .op(n19178) );
  or2_1 U21821 ( .ip1(n19178), .ip2(n19177), .op(n19179) );
  nand2_1 U21822 ( .ip1(n19180), .ip2(n19179), .op(n19181) );
  xnor2_1 U21823 ( .ip1(n19182), .ip2(n19181), .op(n19183) );
  nand2_1 U21824 ( .ip1(n19183), .ip2(n21577), .op(n19215) );
  nor3_1 U21825 ( .ip1(n19186), .ip2(n19185), .ip3(n19184), .op(n19211) );
  inv_1 U21826 ( .ip(n20884), .op(n19192) );
  nand4_1 U21827 ( .ip1(n19190), .ip2(n19189), .ip3(n19188), .ip4(n19187), 
        .op(n20886) );
  nor2_1 U21828 ( .ip1(n18918), .ip2(n20886), .op(n19191) );
  not_ab_or_c_or_d U21829 ( .ip1(n20896), .ip2(n19192), .ip3(n19191), .ip4(
        n20724), .op(n19197) );
  nand2_1 U21830 ( .ip1(n19194), .ip2(n19193), .op(n19196) );
  nand2_1 U21831 ( .ip1(n20897), .ip2(n21540), .op(n19195) );
  nand3_1 U21832 ( .ip1(n19197), .ip2(n19196), .ip3(n19195), .op(n19209) );
  inv_1 U21833 ( .ip(n19199), .op(n19198) );
  nor3_1 U21834 ( .ip1(n13743), .ip2(n21551), .ip3(n19198), .op(n19202) );
  nor2_1 U21835 ( .ip1(n13601), .ip2(n19199), .op(n19200) );
  nor2_1 U21836 ( .ip1(n20907), .ip2(n19200), .op(n19201) );
  not_ab_or_c_or_d U21837 ( .ip1(n20911), .ip2(n19203), .ip3(n19202), .ip4(
        n19201), .op(n19207) );
  nand3_1 U21838 ( .ip1(n19205), .ip2(n19204), .ip3(n19427), .op(n19206) );
  nand4_1 U21839 ( .ip1(n19209), .ip2(n19208), .ip3(n19207), .ip4(n19206), 
        .op(n19210) );
  not_ab_or_c_or_d U21840 ( .ip1(n19213), .ip2(n19212), .ip3(n19211), .ip4(
        n19210), .op(n19214) );
  nand2_1 U21841 ( .ip1(n19215), .ip2(n19214), .op(dmem_haddr[27]) );
  mux2_1 U21842 ( .ip1(dmem_haddr[27]), .ip2(\pipeline/alu_out_WB [27]), .s(
        n19505), .op(n8705) );
  inv_1 U21843 ( .ip(n19216), .op(n19217) );
  nor2_1 U21844 ( .ip1(\pipeline/csr/time_full [27]), .ip2(n19217), .op(n19219) );
  nor3_1 U21845 ( .ip1(n21177), .ip2(n19254), .ip3(n19219), .op(n19218) );
  not_ab_or_c_or_d U21846 ( .ip1(n21179), .ip2(n19243), .ip3(n21217), .ip4(
        n19218), .op(n19222) );
  nor2_1 U21847 ( .ip1(n19219), .ip2(n19254), .op(n19220) );
  nor2_1 U21848 ( .ip1(n21198), .ip2(n19220), .op(n19221) );
  nor2_1 U21849 ( .ip1(n19222), .ip2(n19221), .op(\pipeline/csr/N1964 ) );
  inv_1 U21850 ( .ip(n19223), .op(n19224) );
  nor2_1 U21851 ( .ip1(\pipeline/csr/cycle_full [27]), .ip2(n19224), .op(
        n19226) );
  nor3_1 U21852 ( .ip1(n19276), .ip2(n19226), .ip3(n21215), .op(n19225) );
  not_ab_or_c_or_d U21853 ( .ip1(n21076), .ip2(n19243), .ip3(n21120), .ip4(
        n19225), .op(n19229) );
  nor2_1 U21854 ( .ip1(n19226), .ip2(n19276), .op(n19227) );
  nor2_1 U21855 ( .ip1(n21198), .ip2(n19227), .op(n19228) );
  nor2_1 U21856 ( .ip1(n19229), .ip2(n19228), .op(\pipeline/csr/N1900 ) );
  nand2_1 U21857 ( .ip1(\pipeline/csr/mtimecmp [27]), .ip2(n22363), .op(n19231) );
  nand2_1 U21858 ( .ip1(n22365), .ip2(n19243), .op(n19230) );
  nand2_1 U21859 ( .ip1(n19231), .ip2(n19230), .op(n9995) );
  nand2_1 U21860 ( .ip1(\pipeline/csr/mie [27]), .ip2(n22356), .op(n19233) );
  nand2_1 U21861 ( .ip1(n22357), .ip2(n19243), .op(n19232) );
  nand2_1 U21862 ( .ip1(n19233), .ip2(n19232), .op(n10033) );
  inv_1 U21863 ( .ip(n19243), .op(n19234) );
  nor2_1 U21864 ( .ip1(n19234), .ip2(n22305), .op(n19238) );
  not_ab_or_c_or_d U21865 ( .ip1(n19236), .ip2(n19235), .ip3(n19294), .ip4(
        n22308), .op(n19237) );
  or2_1 U21866 ( .ip1(n19238), .ip2(n19237), .op(\pipeline/csr/N1932 ) );
  nand2_1 U21867 ( .ip1(n22282), .ip2(n19243), .op(n19242) );
  xnor2_1 U21868 ( .ip1(\pipeline/csr/time_full [59]), .ip2(n19239), .op(
        n19240) );
  nand2_1 U21869 ( .ip1(n22284), .ip2(n19240), .op(n19241) );
  nand2_1 U21870 ( .ip1(n19242), .ip2(n19241), .op(\pipeline/csr/N1996 ) );
  nand2_1 U21871 ( .ip1(n20844), .ip2(n19243), .op(n19248) );
  nand2_1 U21872 ( .ip1(n21117), .ip2(\pipeline/csr/instret_full [59]), .op(
        n19247) );
  or2_1 U21873 ( .ip1(\pipeline/csr/instret_full [59]), .ip2(n19244), .op(
        n19245) );
  nand3_1 U21874 ( .ip1(n20334), .ip2(n19250), .ip3(n19245), .op(n19246) );
  nand3_1 U21875 ( .ip1(n19248), .ip2(n19247), .ip3(n19246), .op(n10079) );
  nor2_1 U21876 ( .ip1(n22229), .ip2(n21110), .op(n19253) );
  not_ab_or_c_or_d U21877 ( .ip1(n19251), .ip2(n19250), .ip3(n19249), .ip4(
        n21111), .op(n19252) );
  ab_or_c_or_d U21878 ( .ip1(\pipeline/csr/instret_full [60]), .ip2(n21117), 
        .ip3(n19253), .ip4(n19252), .op(n10078) );
  or2_1 U21879 ( .ip1(\pipeline/csr/time_full [28]), .ip2(n19254), .op(n19255)
         );
  nand2_1 U21880 ( .ip1(n19256), .ip2(n19255), .op(n19258) );
  nor2_1 U21881 ( .ip1(n21177), .ip2(n19258), .op(n19257) );
  not_ab_or_c_or_d U21882 ( .ip1(n21179), .ip2(n22281), .ip3(n21120), .ip4(
        n19257), .op(n19261) );
  inv_1 U21883 ( .ip(n19258), .op(n19259) );
  nor2_1 U21884 ( .ip1(n21198), .ip2(n19259), .op(n19260) );
  nor2_1 U21885 ( .ip1(n19261), .ip2(n19260), .op(\pipeline/csr/N1965 ) );
  inv_1 U21886 ( .ip(n19262), .op(n19263) );
  nor2_1 U21887 ( .ip1(\pipeline/csr/mtime_full [28]), .ip2(n19263), .op(
        n19266) );
  nor3_1 U21888 ( .ip1(n21193), .ip2(n19266), .ip3(n19265), .op(n19264) );
  not_ab_or_c_or_d U21889 ( .ip1(n21195), .ip2(n22281), .ip3(n21120), .ip4(
        n19264), .op(n19269) );
  nor2_1 U21890 ( .ip1(n19266), .ip2(n19265), .op(n19267) );
  nor2_1 U21891 ( .ip1(n22254), .ip2(n19267), .op(n19268) );
  nor2_1 U21892 ( .ip1(n19269), .ip2(n19268), .op(\pipeline/csr/N2109 ) );
  nand2_1 U21893 ( .ip1(\pipeline/csr/mscratch [28]), .ip2(n22013), .op(n19271) );
  nand2_1 U21894 ( .ip1(n22014), .ip2(n22281), .op(n19270) );
  nand2_1 U21895 ( .ip1(n19271), .ip2(n19270), .op(n9900) );
  nand2_1 U21896 ( .ip1(\pipeline/csr/from_host [28]), .ip2(n22372), .op(
        n19273) );
  nand2_1 U21897 ( .ip1(n22373), .ip2(n22281), .op(n19272) );
  nand2_1 U21898 ( .ip1(n19273), .ip2(n19272), .op(n9932) );
  nand2_1 U21899 ( .ip1(n22378), .ip2(n22281), .op(n19275) );
  nand2_1 U21900 ( .ip1(\pipeline/csr/to_host [28]), .ip2(n22376), .op(n19274)
         );
  nand2_1 U21901 ( .ip1(n19275), .ip2(n19274), .op(n8744) );
  or2_1 U21902 ( .ip1(\pipeline/csr/cycle_full [28]), .ip2(n19276), .op(n19277) );
  nand2_1 U21903 ( .ip1(n19278), .ip2(n19277), .op(n19279) );
  or2_1 U21904 ( .ip1(n21145), .ip2(n19279), .op(n19281) );
  nand2_1 U21905 ( .ip1(n22021), .ip2(n22281), .op(n19280) );
  nand2_1 U21906 ( .ip1(n19281), .ip2(n19280), .op(\pipeline/csr/N1901 ) );
  nand2_1 U21907 ( .ip1(\pipeline/csr/mtimecmp [28]), .ip2(n22363), .op(n19283) );
  nand2_1 U21908 ( .ip1(n22365), .ip2(n22281), .op(n19282) );
  nand2_1 U21909 ( .ip1(n19283), .ip2(n19282), .op(n9994) );
  mux2_1 U21910 ( .ip1(\pipeline/csr/instret_full [28]), .ip2(n19287), .s(
        n19284), .op(n19286) );
  nor2_1 U21911 ( .ip1(n21012), .ip2(n21011), .op(n19285) );
  nor2_1 U21912 ( .ip1(n19286), .ip2(n19285), .op(n19289) );
  nor2_1 U21913 ( .ip1(n19287), .ip2(n20990), .op(n19288) );
  nor2_1 U21914 ( .ip1(n19289), .ip2(n19288), .op(n19291) );
  nand2_1 U21915 ( .ip1(n21019), .ip2(n22281), .op(n19290) );
  nand2_1 U21916 ( .ip1(n19291), .ip2(n19290), .op(n10110) );
  nand2_1 U21917 ( .ip1(\pipeline/csr/mie [28]), .ip2(n22356), .op(n19293) );
  nand2_1 U21918 ( .ip1(n22357), .ip2(n22281), .op(n19292) );
  nand2_1 U21919 ( .ip1(n19293), .ip2(n19292), .op(n10032) );
  nand2_1 U21920 ( .ip1(n22314), .ip2(n22281), .op(n19298) );
  or2_1 U21921 ( .ip1(\pipeline/csr/cycle_full [60]), .ip2(n19294), .op(n19295) );
  nand3_1 U21922 ( .ip1(n19296), .ip2(n19295), .ip3(n22316), .op(n19297) );
  nand2_1 U21923 ( .ip1(n19298), .ip2(n19297), .op(\pipeline/csr/N1933 ) );
  inv_1 U21924 ( .ip(n19299), .op(n19300) );
  mux2_1 U21925 ( .ip1(\pipeline/csr_rdata_WB [28]), .ip2(n19300), .s(n17429), 
        .op(n8778) );
  nand2_1 U21926 ( .ip1(n19301), .ip2(n21583), .op(n19306) );
  inv_1 U21927 ( .ip(n19302), .op(n19304) );
  nand2_1 U21928 ( .ip1(n19304), .ip2(n19303), .op(n19305) );
  nand3_1 U21929 ( .ip1(n21588), .ip2(n19306), .ip3(n19305), .op(n19307) );
  mux2_1 U21930 ( .ip1(\pipeline/regfile/data[29][23] ), .ip2(n19307), .s(
        n19353), .op(n8977) );
  mux2_1 U21931 ( .ip1(\pipeline/regfile/data[14][23] ), .ip2(n19307), .s(
        n19354), .op(n9457) );
  mux2_1 U21932 ( .ip1(\pipeline/regfile/data[22][23] ), .ip2(n19307), .s(
        n19355), .op(n9201) );
  mux2_1 U21933 ( .ip1(\pipeline/regfile/data[5][23] ), .ip2(n19307), .s(
        n19356), .op(n9745) );
  mux2_1 U21934 ( .ip1(\pipeline/regfile/data[27][23] ), .ip2(n19307), .s(
        n19357), .op(n9041) );
  mux2_1 U21935 ( .ip1(\pipeline/regfile/data[26][23] ), .ip2(n19307), .s(
        n19358), .op(n9073) );
  mux2_1 U21936 ( .ip1(\pipeline/regfile/data[28][23] ), .ip2(n19307), .s(
        n19359), .op(n9009) );
  mux2_1 U21937 ( .ip1(\pipeline/regfile/data[31][23] ), .ip2(n19307), .s(
        n19360), .op(n8913) );
  mux2_1 U21938 ( .ip1(\pipeline/regfile/data[19][23] ), .ip2(n19307), .s(
        n19361), .op(n9297) );
  mux2_1 U21939 ( .ip1(\pipeline/regfile/data[6][23] ), .ip2(n19307), .s(
        n19362), .op(n9713) );
  mux2_1 U21940 ( .ip1(\pipeline/regfile/data[30][23] ), .ip2(n19307), .s(
        n19363), .op(n8945) );
  mux2_1 U21941 ( .ip1(\pipeline/regfile/data[18][23] ), .ip2(n19307), .s(
        n19364), .op(n9329) );
  mux2_1 U21942 ( .ip1(\pipeline/regfile/data[11][23] ), .ip2(n19307), .s(
        n19365), .op(n9553) );
  mux2_1 U21943 ( .ip1(\pipeline/regfile/data[25][23] ), .ip2(n19307), .s(
        n19366), .op(n9105) );
  mux2_1 U21944 ( .ip1(\pipeline/regfile/data[13][23] ), .ip2(n19307), .s(
        n19367), .op(n9489) );
  mux2_1 U21945 ( .ip1(\pipeline/regfile/data[17][23] ), .ip2(n19307), .s(
        n19368), .op(n9361) );
  mux2_1 U21946 ( .ip1(\pipeline/regfile/data[23][23] ), .ip2(n19307), .s(
        n19369), .op(n9169) );
  mux2_1 U21947 ( .ip1(\pipeline/regfile/data[12][23] ), .ip2(n19307), .s(
        n19370), .op(n9521) );
  mux2_1 U21948 ( .ip1(\pipeline/regfile/data[7][23] ), .ip2(n19307), .s(
        n19371), .op(n9681) );
  mux2_1 U21949 ( .ip1(\pipeline/regfile/data[8][23] ), .ip2(n19307), .s(
        n19372), .op(n9649) );
  mux2_1 U21950 ( .ip1(\pipeline/regfile/data[15][23] ), .ip2(n19307), .s(
        n19373), .op(n9425) );
  mux2_1 U21951 ( .ip1(\pipeline/regfile/data[10][23] ), .ip2(n19307), .s(
        n19374), .op(n9585) );
  mux2_1 U21952 ( .ip1(\pipeline/regfile/data[21][23] ), .ip2(n19307), .s(
        n19375), .op(n9233) );
  mux2_1 U21953 ( .ip1(\pipeline/regfile/data[24][23] ), .ip2(n19307), .s(
        n19376), .op(n9137) );
  mux2_1 U21954 ( .ip1(\pipeline/regfile/data[20][23] ), .ip2(n19307), .s(
        n19377), .op(n9265) );
  mux2_1 U21955 ( .ip1(\pipeline/regfile/data[9][23] ), .ip2(n19307), .s(
        n19378), .op(n9617) );
  mux2_1 U21956 ( .ip1(\pipeline/regfile/data[16][23] ), .ip2(n19307), .s(
        n19379), .op(n9393) );
  mux2_1 U21957 ( .ip1(\pipeline/regfile/data[3][23] ), .ip2(n19307), .s(
        n19380), .op(n9809) );
  mux2_1 U21958 ( .ip1(\pipeline/regfile/data[1][23] ), .ip2(n19307), .s(
        n19381), .op(n9873) );
  mux2_1 U21959 ( .ip1(\pipeline/regfile/data[2][23] ), .ip2(n19307), .s(
        n19382), .op(n9841) );
  mux2_1 U21960 ( .ip1(\pipeline/regfile/data[4][23] ), .ip2(n19307), .s(
        n19383), .op(n9777) );
  nand2_1 U21961 ( .ip1(dmem_rdata[22]), .ip2(n21585), .op(n19311) );
  nand2_1 U21962 ( .ip1(n19308), .ip2(n21583), .op(n19310) );
  nand2_1 U21963 ( .ip1(dmem_rdata[30]), .ip2(n19324), .op(n19309) );
  nand4_1 U21964 ( .ip1(n21588), .ip2(n19311), .ip3(n19310), .ip4(n19309), 
        .op(n19312) );
  mux2_1 U21965 ( .ip1(\pipeline/regfile/data[29][22] ), .ip2(n19312), .s(
        n19353), .op(n8978) );
  mux2_1 U21966 ( .ip1(\pipeline/regfile/data[14][22] ), .ip2(n19312), .s(
        n19354), .op(n9458) );
  mux2_1 U21967 ( .ip1(\pipeline/regfile/data[22][22] ), .ip2(n19312), .s(
        n19355), .op(n9202) );
  mux2_1 U21968 ( .ip1(\pipeline/regfile/data[5][22] ), .ip2(n19312), .s(
        n19356), .op(n9746) );
  mux2_1 U21969 ( .ip1(\pipeline/regfile/data[27][22] ), .ip2(n19312), .s(
        n19357), .op(n9042) );
  mux2_1 U21970 ( .ip1(\pipeline/regfile/data[26][22] ), .ip2(n19312), .s(
        n19358), .op(n9074) );
  mux2_1 U21971 ( .ip1(\pipeline/regfile/data[28][22] ), .ip2(n19312), .s(
        n19359), .op(n9010) );
  mux2_1 U21972 ( .ip1(\pipeline/regfile/data[31][22] ), .ip2(n19312), .s(
        n19360), .op(n8914) );
  mux2_1 U21973 ( .ip1(\pipeline/regfile/data[19][22] ), .ip2(n19312), .s(
        n19361), .op(n9298) );
  mux2_1 U21974 ( .ip1(\pipeline/regfile/data[6][22] ), .ip2(n19312), .s(
        n19362), .op(n9714) );
  mux2_1 U21975 ( .ip1(\pipeline/regfile/data[30][22] ), .ip2(n19312), .s(
        n19363), .op(n8946) );
  mux2_1 U21976 ( .ip1(\pipeline/regfile/data[18][22] ), .ip2(n19312), .s(
        n19364), .op(n9330) );
  mux2_1 U21977 ( .ip1(\pipeline/regfile/data[11][22] ), .ip2(n19312), .s(
        n19365), .op(n9554) );
  mux2_1 U21978 ( .ip1(\pipeline/regfile/data[25][22] ), .ip2(n19312), .s(
        n19366), .op(n9106) );
  mux2_1 U21979 ( .ip1(\pipeline/regfile/data[13][22] ), .ip2(n19312), .s(
        n19367), .op(n9490) );
  mux2_1 U21980 ( .ip1(\pipeline/regfile/data[17][22] ), .ip2(n19312), .s(
        n19368), .op(n9362) );
  mux2_1 U21981 ( .ip1(\pipeline/regfile/data[23][22] ), .ip2(n19312), .s(
        n19369), .op(n9170) );
  mux2_1 U21982 ( .ip1(\pipeline/regfile/data[12][22] ), .ip2(n19312), .s(
        n19370), .op(n9522) );
  mux2_1 U21983 ( .ip1(\pipeline/regfile/data[7][22] ), .ip2(n19312), .s(
        n19371), .op(n9682) );
  mux2_1 U21984 ( .ip1(\pipeline/regfile/data[8][22] ), .ip2(n19312), .s(
        n19372), .op(n9650) );
  mux2_1 U21985 ( .ip1(\pipeline/regfile/data[15][22] ), .ip2(n19312), .s(
        n19373), .op(n9426) );
  mux2_1 U21986 ( .ip1(\pipeline/regfile/data[10][22] ), .ip2(n19312), .s(
        n19374), .op(n9586) );
  mux2_1 U21987 ( .ip1(\pipeline/regfile/data[21][22] ), .ip2(n19312), .s(
        n19375), .op(n9234) );
  mux2_1 U21988 ( .ip1(\pipeline/regfile/data[24][22] ), .ip2(n19312), .s(
        n19376), .op(n9138) );
  mux2_1 U21989 ( .ip1(\pipeline/regfile/data[20][22] ), .ip2(n19312), .s(
        n19377), .op(n9266) );
  mux2_1 U21990 ( .ip1(\pipeline/regfile/data[9][22] ), .ip2(n19312), .s(
        n19378), .op(n9618) );
  mux2_1 U21991 ( .ip1(\pipeline/regfile/data[16][22] ), .ip2(n19312), .s(
        n19379), .op(n9394) );
  mux2_1 U21992 ( .ip1(\pipeline/regfile/data[3][22] ), .ip2(n19312), .s(
        n19380), .op(n9810) );
  mux2_1 U21993 ( .ip1(\pipeline/regfile/data[1][22] ), .ip2(n19312), .s(
        n19381), .op(n9874) );
  mux2_1 U21994 ( .ip1(\pipeline/regfile/data[2][22] ), .ip2(n19312), .s(
        n19382), .op(n9842) );
  mux2_1 U21995 ( .ip1(\pipeline/regfile/data[4][22] ), .ip2(n19312), .s(
        n19383), .op(n9778) );
  nand2_1 U21996 ( .ip1(dmem_rdata[20]), .ip2(n21585), .op(n19316) );
  nand2_1 U21997 ( .ip1(n19313), .ip2(n21583), .op(n19315) );
  nand2_1 U21998 ( .ip1(dmem_rdata[28]), .ip2(n19324), .op(n19314) );
  nand4_1 U21999 ( .ip1(n21588), .ip2(n19316), .ip3(n19315), .ip4(n19314), 
        .op(n19317) );
  mux2_1 U22000 ( .ip1(\pipeline/regfile/data[29][20] ), .ip2(n19317), .s(
        n19353), .op(n8980) );
  mux2_1 U22001 ( .ip1(\pipeline/regfile/data[14][20] ), .ip2(n19317), .s(
        n19354), .op(n9460) );
  mux2_1 U22002 ( .ip1(\pipeline/regfile/data[22][20] ), .ip2(n19317), .s(
        n19355), .op(n9204) );
  mux2_1 U22003 ( .ip1(\pipeline/regfile/data[5][20] ), .ip2(n19317), .s(
        n19356), .op(n9748) );
  mux2_1 U22004 ( .ip1(\pipeline/regfile/data[27][20] ), .ip2(n19317), .s(
        n19357), .op(n9044) );
  mux2_1 U22005 ( .ip1(\pipeline/regfile/data[26][20] ), .ip2(n19317), .s(
        n19358), .op(n9076) );
  mux2_1 U22006 ( .ip1(\pipeline/regfile/data[28][20] ), .ip2(n19317), .s(
        n19359), .op(n9012) );
  mux2_1 U22007 ( .ip1(\pipeline/regfile/data[31][20] ), .ip2(n19317), .s(
        n19360), .op(n8916) );
  mux2_1 U22008 ( .ip1(\pipeline/regfile/data[19][20] ), .ip2(n19317), .s(
        n19361), .op(n9300) );
  mux2_1 U22009 ( .ip1(\pipeline/regfile/data[6][20] ), .ip2(n19317), .s(
        n19362), .op(n9716) );
  mux2_1 U22010 ( .ip1(\pipeline/regfile/data[30][20] ), .ip2(n19317), .s(
        n19363), .op(n8948) );
  mux2_1 U22011 ( .ip1(\pipeline/regfile/data[18][20] ), .ip2(n19317), .s(
        n19364), .op(n9332) );
  mux2_1 U22012 ( .ip1(\pipeline/regfile/data[11][20] ), .ip2(n19317), .s(
        n19365), .op(n9556) );
  mux2_1 U22013 ( .ip1(\pipeline/regfile/data[25][20] ), .ip2(n19317), .s(
        n19366), .op(n9108) );
  mux2_1 U22014 ( .ip1(\pipeline/regfile/data[13][20] ), .ip2(n19317), .s(
        n19367), .op(n9492) );
  mux2_1 U22015 ( .ip1(\pipeline/regfile/data[17][20] ), .ip2(n19317), .s(
        n19368), .op(n9364) );
  mux2_1 U22016 ( .ip1(\pipeline/regfile/data[23][20] ), .ip2(n19317), .s(
        n19369), .op(n9172) );
  mux2_1 U22017 ( .ip1(\pipeline/regfile/data[12][20] ), .ip2(n19317), .s(
        n19370), .op(n9524) );
  mux2_1 U22018 ( .ip1(\pipeline/regfile/data[7][20] ), .ip2(n19317), .s(
        n19371), .op(n9684) );
  mux2_1 U22019 ( .ip1(\pipeline/regfile/data[8][20] ), .ip2(n19317), .s(
        n19372), .op(n9652) );
  mux2_1 U22020 ( .ip1(\pipeline/regfile/data[15][20] ), .ip2(n19317), .s(
        n19373), .op(n9428) );
  mux2_1 U22021 ( .ip1(\pipeline/regfile/data[10][20] ), .ip2(n19317), .s(
        n19374), .op(n9588) );
  mux2_1 U22022 ( .ip1(\pipeline/regfile/data[21][20] ), .ip2(n19317), .s(
        n19375), .op(n9236) );
  mux2_1 U22023 ( .ip1(\pipeline/regfile/data[24][20] ), .ip2(n19317), .s(
        n19376), .op(n9140) );
  mux2_1 U22024 ( .ip1(\pipeline/regfile/data[20][20] ), .ip2(n19317), .s(
        n19377), .op(n9268) );
  mux2_1 U22025 ( .ip1(\pipeline/regfile/data[9][20] ), .ip2(n19317), .s(
        n19378), .op(n9620) );
  mux2_1 U22026 ( .ip1(\pipeline/regfile/data[16][20] ), .ip2(n19317), .s(
        n19379), .op(n9396) );
  mux2_1 U22027 ( .ip1(\pipeline/regfile/data[3][20] ), .ip2(n19317), .s(
        n19380), .op(n9812) );
  mux2_1 U22028 ( .ip1(\pipeline/regfile/data[1][20] ), .ip2(n19317), .s(
        n19381), .op(n9876) );
  mux2_1 U22029 ( .ip1(\pipeline/regfile/data[2][20] ), .ip2(n19317), .s(
        n19382), .op(n9844) );
  mux2_1 U22030 ( .ip1(\pipeline/regfile/data[4][20] ), .ip2(n19317), .s(
        n19383), .op(n9780) );
  nand2_1 U22031 ( .ip1(dmem_rdata[17]), .ip2(n21585), .op(n19321) );
  nand2_1 U22032 ( .ip1(n19318), .ip2(n21583), .op(n19320) );
  nand2_1 U22033 ( .ip1(dmem_rdata[25]), .ip2(n19324), .op(n19319) );
  nand4_1 U22034 ( .ip1(n21588), .ip2(n19321), .ip3(n19320), .ip4(n19319), 
        .op(n19322) );
  mux2_1 U22035 ( .ip1(\pipeline/regfile/data[29][17] ), .ip2(n19322), .s(
        n19353), .op(n8983) );
  mux2_1 U22036 ( .ip1(\pipeline/regfile/data[14][17] ), .ip2(n19322), .s(
        n19354), .op(n9463) );
  mux2_1 U22037 ( .ip1(\pipeline/regfile/data[22][17] ), .ip2(n19322), .s(
        n19355), .op(n9207) );
  mux2_1 U22038 ( .ip1(\pipeline/regfile/data[5][17] ), .ip2(n19322), .s(
        n19356), .op(n9751) );
  mux2_1 U22039 ( .ip1(\pipeline/regfile/data[27][17] ), .ip2(n19322), .s(
        n19357), .op(n9047) );
  mux2_1 U22040 ( .ip1(\pipeline/regfile/data[26][17] ), .ip2(n19322), .s(
        n19358), .op(n9079) );
  mux2_1 U22041 ( .ip1(\pipeline/regfile/data[28][17] ), .ip2(n19322), .s(
        n19359), .op(n9015) );
  mux2_1 U22042 ( .ip1(\pipeline/regfile/data[31][17] ), .ip2(n19322), .s(
        n19360), .op(n8919) );
  mux2_1 U22043 ( .ip1(\pipeline/regfile/data[19][17] ), .ip2(n19322), .s(
        n19361), .op(n9303) );
  mux2_1 U22044 ( .ip1(\pipeline/regfile/data[6][17] ), .ip2(n19322), .s(
        n19362), .op(n9719) );
  mux2_1 U22045 ( .ip1(\pipeline/regfile/data[30][17] ), .ip2(n19322), .s(
        n19363), .op(n8951) );
  mux2_1 U22046 ( .ip1(\pipeline/regfile/data[18][17] ), .ip2(n19322), .s(
        n19364), .op(n9335) );
  mux2_1 U22047 ( .ip1(\pipeline/regfile/data[11][17] ), .ip2(n19322), .s(
        n19365), .op(n9559) );
  mux2_1 U22048 ( .ip1(\pipeline/regfile/data[25][17] ), .ip2(n19322), .s(
        n19366), .op(n9111) );
  mux2_1 U22049 ( .ip1(\pipeline/regfile/data[13][17] ), .ip2(n19322), .s(
        n19367), .op(n9495) );
  mux2_1 U22050 ( .ip1(\pipeline/regfile/data[17][17] ), .ip2(n19322), .s(
        n19368), .op(n9367) );
  mux2_1 U22051 ( .ip1(\pipeline/regfile/data[23][17] ), .ip2(n19322), .s(
        n19369), .op(n9175) );
  mux2_1 U22052 ( .ip1(\pipeline/regfile/data[12][17] ), .ip2(n19322), .s(
        n19370), .op(n9527) );
  mux2_1 U22053 ( .ip1(\pipeline/regfile/data[7][17] ), .ip2(n19322), .s(
        n19371), .op(n9687) );
  mux2_1 U22054 ( .ip1(\pipeline/regfile/data[8][17] ), .ip2(n19322), .s(
        n19372), .op(n9655) );
  mux2_1 U22055 ( .ip1(\pipeline/regfile/data[15][17] ), .ip2(n19322), .s(
        n19373), .op(n9431) );
  mux2_1 U22056 ( .ip1(\pipeline/regfile/data[10][17] ), .ip2(n19322), .s(
        n19374), .op(n9591) );
  mux2_1 U22057 ( .ip1(\pipeline/regfile/data[21][17] ), .ip2(n19322), .s(
        n19375), .op(n9239) );
  mux2_1 U22058 ( .ip1(\pipeline/regfile/data[24][17] ), .ip2(n19322), .s(
        n19376), .op(n9143) );
  mux2_1 U22059 ( .ip1(\pipeline/regfile/data[20][17] ), .ip2(n19322), .s(
        n19377), .op(n9271) );
  mux2_1 U22060 ( .ip1(\pipeline/regfile/data[9][17] ), .ip2(n19322), .s(
        n19378), .op(n9623) );
  mux2_1 U22061 ( .ip1(\pipeline/regfile/data[16][17] ), .ip2(n19322), .s(
        n19379), .op(n9399) );
  mux2_1 U22062 ( .ip1(\pipeline/regfile/data[3][17] ), .ip2(n19322), .s(
        n19380), .op(n9815) );
  mux2_1 U22063 ( .ip1(\pipeline/regfile/data[1][17] ), .ip2(n19322), .s(
        n19381), .op(n9879) );
  mux2_1 U22064 ( .ip1(\pipeline/regfile/data[2][17] ), .ip2(n19322), .s(
        n19382), .op(n9847) );
  mux2_1 U22065 ( .ip1(\pipeline/regfile/data[4][17] ), .ip2(n19322), .s(
        n19383), .op(n9783) );
  nand2_1 U22066 ( .ip1(n21585), .ip2(dmem_rdata[16]), .op(n19327) );
  nand2_1 U22067 ( .ip1(n19323), .ip2(n21583), .op(n19326) );
  nand2_1 U22068 ( .ip1(n19324), .ip2(dmem_rdata[24]), .op(n19325) );
  nand4_1 U22069 ( .ip1(n21588), .ip2(n19327), .ip3(n19326), .ip4(n19325), 
        .op(n19328) );
  mux2_1 U22070 ( .ip1(\pipeline/regfile/data[29][16] ), .ip2(n19328), .s(
        n19353), .op(n8984) );
  mux2_1 U22071 ( .ip1(\pipeline/regfile/data[14][16] ), .ip2(n19328), .s(
        n19354), .op(n9464) );
  mux2_1 U22072 ( .ip1(\pipeline/regfile/data[22][16] ), .ip2(n19328), .s(
        n19355), .op(n9208) );
  mux2_1 U22073 ( .ip1(\pipeline/regfile/data[5][16] ), .ip2(n19328), .s(
        n19356), .op(n9752) );
  mux2_1 U22074 ( .ip1(\pipeline/regfile/data[27][16] ), .ip2(n19328), .s(
        n19357), .op(n9048) );
  mux2_1 U22075 ( .ip1(\pipeline/regfile/data[26][16] ), .ip2(n19328), .s(
        n19358), .op(n9080) );
  mux2_1 U22076 ( .ip1(\pipeline/regfile/data[28][16] ), .ip2(n19328), .s(
        n19359), .op(n9016) );
  mux2_1 U22077 ( .ip1(\pipeline/regfile/data[31][16] ), .ip2(n19328), .s(
        n19360), .op(n8920) );
  mux2_1 U22078 ( .ip1(\pipeline/regfile/data[19][16] ), .ip2(n19328), .s(
        n19361), .op(n9304) );
  mux2_1 U22079 ( .ip1(\pipeline/regfile/data[6][16] ), .ip2(n19328), .s(
        n19362), .op(n9720) );
  mux2_1 U22080 ( .ip1(\pipeline/regfile/data[30][16] ), .ip2(n19328), .s(
        n19363), .op(n8952) );
  mux2_1 U22081 ( .ip1(\pipeline/regfile/data[18][16] ), .ip2(n19328), .s(
        n19364), .op(n9336) );
  mux2_1 U22082 ( .ip1(\pipeline/regfile/data[11][16] ), .ip2(n19328), .s(
        n19365), .op(n9560) );
  mux2_1 U22083 ( .ip1(\pipeline/regfile/data[25][16] ), .ip2(n19328), .s(
        n19366), .op(n9112) );
  mux2_1 U22084 ( .ip1(\pipeline/regfile/data[13][16] ), .ip2(n19328), .s(
        n19367), .op(n9496) );
  mux2_1 U22085 ( .ip1(\pipeline/regfile/data[17][16] ), .ip2(n19328), .s(
        n19368), .op(n9368) );
  mux2_1 U22086 ( .ip1(\pipeline/regfile/data[23][16] ), .ip2(n19328), .s(
        n19369), .op(n9176) );
  mux2_1 U22087 ( .ip1(\pipeline/regfile/data[12][16] ), .ip2(n19328), .s(
        n19370), .op(n9528) );
  mux2_1 U22088 ( .ip1(\pipeline/regfile/data[7][16] ), .ip2(n19328), .s(
        n19371), .op(n9688) );
  mux2_1 U22089 ( .ip1(\pipeline/regfile/data[8][16] ), .ip2(n19328), .s(
        n19372), .op(n9656) );
  mux2_1 U22090 ( .ip1(\pipeline/regfile/data[15][16] ), .ip2(n19328), .s(
        n19373), .op(n9432) );
  mux2_1 U22091 ( .ip1(\pipeline/regfile/data[10][16] ), .ip2(n19328), .s(
        n19374), .op(n9592) );
  mux2_1 U22092 ( .ip1(\pipeline/regfile/data[21][16] ), .ip2(n19328), .s(
        n19375), .op(n9240) );
  mux2_1 U22093 ( .ip1(\pipeline/regfile/data[24][16] ), .ip2(n19328), .s(
        n19376), .op(n9144) );
  mux2_1 U22094 ( .ip1(\pipeline/regfile/data[20][16] ), .ip2(n19328), .s(
        n19377), .op(n9272) );
  mux2_1 U22095 ( .ip1(\pipeline/regfile/data[9][16] ), .ip2(n19328), .s(
        n19378), .op(n9624) );
  mux2_1 U22096 ( .ip1(\pipeline/regfile/data[16][16] ), .ip2(n19328), .s(
        n19379), .op(n9400) );
  mux2_1 U22097 ( .ip1(\pipeline/regfile/data[3][16] ), .ip2(n19328), .s(
        n19380), .op(n9816) );
  mux2_1 U22098 ( .ip1(\pipeline/regfile/data[1][16] ), .ip2(n19328), .s(
        n19381), .op(n9880) );
  mux2_1 U22099 ( .ip1(\pipeline/regfile/data[2][16] ), .ip2(n19328), .s(
        n19382), .op(n9848) );
  mux2_1 U22100 ( .ip1(\pipeline/regfile/data[4][16] ), .ip2(n19328), .s(
        n19383), .op(n9784) );
  nor2_1 U22101 ( .ip1(n22071), .ip2(n21235), .op(n19409) );
  nand2_1 U22102 ( .ip1(n21238), .ip2(dmem_rdata[14]), .op(n19329) );
  nor2_1 U22103 ( .ip1(n22071), .ip2(n19329), .op(n19333) );
  inv_1 U22104 ( .ip(n19330), .op(n19331) );
  nor2_1 U22105 ( .ip1(n19331), .ip2(n19404), .op(n19332) );
  not_ab_or_c_or_d U22106 ( .ip1(dmem_rdata[22]), .ip2(n19409), .ip3(n19333), 
        .ip4(n19332), .op(n19335) );
  inv_1 U22107 ( .ip(n19390), .op(n19412) );
  nand2_1 U22108 ( .ip1(dmem_rdata[30]), .ip2(n19410), .op(n19334) );
  nand3_1 U22109 ( .ip1(n19335), .ip2(n19412), .ip3(n19334), .op(n19336) );
  mux2_1 U22110 ( .ip1(\pipeline/regfile/data[29][14] ), .ip2(n19336), .s(
        n19353), .op(n8986) );
  mux2_1 U22111 ( .ip1(\pipeline/regfile/data[14][14] ), .ip2(n19336), .s(
        n19354), .op(n9466) );
  mux2_1 U22112 ( .ip1(\pipeline/regfile/data[22][14] ), .ip2(n19336), .s(
        n19355), .op(n9210) );
  mux2_1 U22113 ( .ip1(\pipeline/regfile/data[5][14] ), .ip2(n19336), .s(
        n19356), .op(n9754) );
  mux2_1 U22114 ( .ip1(\pipeline/regfile/data[27][14] ), .ip2(n19336), .s(
        n19357), .op(n9050) );
  mux2_1 U22115 ( .ip1(\pipeline/regfile/data[26][14] ), .ip2(n19336), .s(
        n19358), .op(n9082) );
  mux2_1 U22116 ( .ip1(\pipeline/regfile/data[28][14] ), .ip2(n19336), .s(
        n19359), .op(n9018) );
  mux2_1 U22117 ( .ip1(\pipeline/regfile/data[31][14] ), .ip2(n19336), .s(
        n19360), .op(n8922) );
  mux2_1 U22118 ( .ip1(\pipeline/regfile/data[19][14] ), .ip2(n19336), .s(
        n19361), .op(n9306) );
  mux2_1 U22119 ( .ip1(\pipeline/regfile/data[6][14] ), .ip2(n19336), .s(
        n19362), .op(n9722) );
  mux2_1 U22120 ( .ip1(\pipeline/regfile/data[30][14] ), .ip2(n19336), .s(
        n19363), .op(n8954) );
  mux2_1 U22121 ( .ip1(\pipeline/regfile/data[18][14] ), .ip2(n19336), .s(
        n19364), .op(n9338) );
  mux2_1 U22122 ( .ip1(\pipeline/regfile/data[11][14] ), .ip2(n19336), .s(
        n19365), .op(n9562) );
  mux2_1 U22123 ( .ip1(\pipeline/regfile/data[25][14] ), .ip2(n19336), .s(
        n19366), .op(n9114) );
  mux2_1 U22124 ( .ip1(\pipeline/regfile/data[13][14] ), .ip2(n19336), .s(
        n19367), .op(n9498) );
  mux2_1 U22125 ( .ip1(\pipeline/regfile/data[17][14] ), .ip2(n19336), .s(
        n19368), .op(n9370) );
  mux2_1 U22126 ( .ip1(\pipeline/regfile/data[23][14] ), .ip2(n19336), .s(
        n19369), .op(n9178) );
  mux2_1 U22127 ( .ip1(\pipeline/regfile/data[12][14] ), .ip2(n19336), .s(
        n19370), .op(n9530) );
  mux2_1 U22128 ( .ip1(\pipeline/regfile/data[7][14] ), .ip2(n19336), .s(
        n19371), .op(n9690) );
  mux2_1 U22129 ( .ip1(\pipeline/regfile/data[8][14] ), .ip2(n19336), .s(
        n19372), .op(n9658) );
  mux2_1 U22130 ( .ip1(\pipeline/regfile/data[15][14] ), .ip2(n19336), .s(
        n19373), .op(n9434) );
  mux2_1 U22131 ( .ip1(\pipeline/regfile/data[10][14] ), .ip2(n19336), .s(
        n19374), .op(n9594) );
  mux2_1 U22132 ( .ip1(\pipeline/regfile/data[21][14] ), .ip2(n19336), .s(
        n19375), .op(n9242) );
  mux2_1 U22133 ( .ip1(\pipeline/regfile/data[24][14] ), .ip2(n19336), .s(
        n19376), .op(n9146) );
  mux2_1 U22134 ( .ip1(\pipeline/regfile/data[20][14] ), .ip2(n19336), .s(
        n19377), .op(n9274) );
  mux2_1 U22135 ( .ip1(\pipeline/regfile/data[9][14] ), .ip2(n19336), .s(
        n19378), .op(n9626) );
  mux2_1 U22136 ( .ip1(\pipeline/regfile/data[16][14] ), .ip2(n19336), .s(
        n19379), .op(n9402) );
  mux2_1 U22137 ( .ip1(\pipeline/regfile/data[3][14] ), .ip2(n19336), .s(
        n19380), .op(n9818) );
  mux2_1 U22138 ( .ip1(\pipeline/regfile/data[1][14] ), .ip2(n19336), .s(
        n19381), .op(n9882) );
  mux2_1 U22139 ( .ip1(\pipeline/regfile/data[2][14] ), .ip2(n19336), .s(
        n19382), .op(n9850) );
  mux2_1 U22140 ( .ip1(\pipeline/regfile/data[4][14] ), .ip2(n19336), .s(
        n19383), .op(n9786) );
  nand2_1 U22141 ( .ip1(n21238), .ip2(dmem_rdata[13]), .op(n19337) );
  or2_1 U22142 ( .ip1(n19337), .ip2(n22071), .op(n19340) );
  nand2_1 U22143 ( .ip1(n19386), .ip2(dmem_rdata[21]), .op(n19338) );
  or2_1 U22144 ( .ip1(n19338), .ip2(n22071), .op(n19339) );
  nand2_1 U22145 ( .ip1(n19340), .ip2(n19339), .op(n19341) );
  not_ab_or_c_or_d U22146 ( .ip1(n19342), .ip2(n21583), .ip3(n19341), .ip4(
        n19390), .op(n19344) );
  nand2_1 U22147 ( .ip1(dmem_rdata[29]), .ip2(n19410), .op(n19343) );
  nand2_1 U22148 ( .ip1(n19344), .ip2(n19343), .op(n19345) );
  mux2_1 U22149 ( .ip1(\pipeline/regfile/data[29][13] ), .ip2(n19345), .s(
        n19353), .op(n8987) );
  mux2_1 U22150 ( .ip1(\pipeline/regfile/data[14][13] ), .ip2(n19345), .s(
        n19354), .op(n9467) );
  mux2_1 U22151 ( .ip1(\pipeline/regfile/data[22][13] ), .ip2(n19345), .s(
        n19355), .op(n9211) );
  mux2_1 U22152 ( .ip1(\pipeline/regfile/data[5][13] ), .ip2(n19345), .s(
        n19356), .op(n9755) );
  mux2_1 U22153 ( .ip1(\pipeline/regfile/data[27][13] ), .ip2(n19345), .s(
        n19357), .op(n9051) );
  mux2_1 U22154 ( .ip1(\pipeline/regfile/data[26][13] ), .ip2(n19345), .s(
        n19358), .op(n9083) );
  mux2_1 U22155 ( .ip1(\pipeline/regfile/data[28][13] ), .ip2(n19345), .s(
        n19359), .op(n9019) );
  mux2_1 U22156 ( .ip1(\pipeline/regfile/data[31][13] ), .ip2(n19345), .s(
        n19360), .op(n8923) );
  mux2_1 U22157 ( .ip1(\pipeline/regfile/data[19][13] ), .ip2(n19345), .s(
        n19361), .op(n9307) );
  mux2_1 U22158 ( .ip1(\pipeline/regfile/data[6][13] ), .ip2(n19345), .s(
        n19362), .op(n9723) );
  mux2_1 U22159 ( .ip1(\pipeline/regfile/data[30][13] ), .ip2(n19345), .s(
        n19363), .op(n8955) );
  mux2_1 U22160 ( .ip1(\pipeline/regfile/data[18][13] ), .ip2(n19345), .s(
        n19364), .op(n9339) );
  mux2_1 U22161 ( .ip1(\pipeline/regfile/data[11][13] ), .ip2(n19345), .s(
        n19365), .op(n9563) );
  mux2_1 U22162 ( .ip1(\pipeline/regfile/data[25][13] ), .ip2(n19345), .s(
        n19366), .op(n9115) );
  mux2_1 U22163 ( .ip1(\pipeline/regfile/data[13][13] ), .ip2(n19345), .s(
        n19367), .op(n9499) );
  mux2_1 U22164 ( .ip1(\pipeline/regfile/data[17][13] ), .ip2(n19345), .s(
        n19368), .op(n9371) );
  mux2_1 U22165 ( .ip1(\pipeline/regfile/data[23][13] ), .ip2(n19345), .s(
        n19369), .op(n9179) );
  mux2_1 U22166 ( .ip1(\pipeline/regfile/data[12][13] ), .ip2(n19345), .s(
        n19370), .op(n9531) );
  mux2_1 U22167 ( .ip1(\pipeline/regfile/data[7][13] ), .ip2(n19345), .s(
        n19371), .op(n9691) );
  mux2_1 U22168 ( .ip1(\pipeline/regfile/data[8][13] ), .ip2(n19345), .s(
        n19372), .op(n9659) );
  mux2_1 U22169 ( .ip1(\pipeline/regfile/data[15][13] ), .ip2(n19345), .s(
        n19373), .op(n9435) );
  mux2_1 U22170 ( .ip1(\pipeline/regfile/data[10][13] ), .ip2(n19345), .s(
        n19374), .op(n9595) );
  mux2_1 U22171 ( .ip1(\pipeline/regfile/data[21][13] ), .ip2(n19345), .s(
        n19375), .op(n9243) );
  mux2_1 U22172 ( .ip1(\pipeline/regfile/data[24][13] ), .ip2(n19345), .s(
        n19376), .op(n9147) );
  mux2_1 U22173 ( .ip1(\pipeline/regfile/data[20][13] ), .ip2(n19345), .s(
        n19377), .op(n9275) );
  mux2_1 U22174 ( .ip1(\pipeline/regfile/data[9][13] ), .ip2(n19345), .s(
        n19378), .op(n9627) );
  mux2_1 U22175 ( .ip1(\pipeline/regfile/data[16][13] ), .ip2(n19345), .s(
        n19379), .op(n9403) );
  mux2_1 U22176 ( .ip1(\pipeline/regfile/data[3][13] ), .ip2(n19345), .s(
        n19380), .op(n9819) );
  mux2_1 U22177 ( .ip1(\pipeline/regfile/data[1][13] ), .ip2(n19345), .s(
        n19381), .op(n9883) );
  mux2_1 U22178 ( .ip1(\pipeline/regfile/data[2][13] ), .ip2(n19345), .s(
        n19382), .op(n9851) );
  mux2_1 U22179 ( .ip1(\pipeline/regfile/data[4][13] ), .ip2(n19345), .s(
        n19383), .op(n9787) );
  inv_1 U22180 ( .ip(n19346), .op(n19347) );
  nor2_1 U22181 ( .ip1(n19347), .ip2(n19404), .op(n19350) );
  nand2_1 U22182 ( .ip1(n21238), .ip2(dmem_rdata[12]), .op(n19348) );
  nor2_1 U22183 ( .ip1(n22071), .ip2(n19348), .op(n19349) );
  not_ab_or_c_or_d U22184 ( .ip1(n19409), .ip2(dmem_rdata[20]), .ip3(n19350), 
        .ip4(n19349), .op(n19352) );
  nand2_1 U22185 ( .ip1(dmem_rdata[28]), .ip2(n19410), .op(n19351) );
  nand3_1 U22186 ( .ip1(n19352), .ip2(n19412), .ip3(n19351), .op(n19384) );
  mux2_1 U22187 ( .ip1(\pipeline/regfile/data[29][12] ), .ip2(n19384), .s(
        n19353), .op(n8988) );
  mux2_1 U22188 ( .ip1(\pipeline/regfile/data[14][12] ), .ip2(n19384), .s(
        n19354), .op(n9468) );
  mux2_1 U22189 ( .ip1(\pipeline/regfile/data[22][12] ), .ip2(n19384), .s(
        n19355), .op(n9212) );
  mux2_1 U22190 ( .ip1(\pipeline/regfile/data[5][12] ), .ip2(n19384), .s(
        n19356), .op(n9756) );
  mux2_1 U22191 ( .ip1(\pipeline/regfile/data[27][12] ), .ip2(n19384), .s(
        n19357), .op(n9052) );
  mux2_1 U22192 ( .ip1(\pipeline/regfile/data[26][12] ), .ip2(n19384), .s(
        n19358), .op(n9084) );
  mux2_1 U22193 ( .ip1(\pipeline/regfile/data[28][12] ), .ip2(n19384), .s(
        n19359), .op(n9020) );
  mux2_1 U22194 ( .ip1(\pipeline/regfile/data[31][12] ), .ip2(n19384), .s(
        n19360), .op(n8924) );
  mux2_1 U22195 ( .ip1(\pipeline/regfile/data[19][12] ), .ip2(n19384), .s(
        n19361), .op(n9308) );
  mux2_1 U22196 ( .ip1(\pipeline/regfile/data[6][12] ), .ip2(n19384), .s(
        n19362), .op(n9724) );
  mux2_1 U22197 ( .ip1(\pipeline/regfile/data[30][12] ), .ip2(n19384), .s(
        n19363), .op(n8956) );
  mux2_1 U22198 ( .ip1(\pipeline/regfile/data[18][12] ), .ip2(n19384), .s(
        n19364), .op(n9340) );
  mux2_1 U22199 ( .ip1(\pipeline/regfile/data[11][12] ), .ip2(n19384), .s(
        n19365), .op(n9564) );
  mux2_1 U22200 ( .ip1(\pipeline/regfile/data[25][12] ), .ip2(n19384), .s(
        n19366), .op(n9116) );
  mux2_1 U22201 ( .ip1(\pipeline/regfile/data[13][12] ), .ip2(n19384), .s(
        n19367), .op(n9500) );
  mux2_1 U22202 ( .ip1(\pipeline/regfile/data[17][12] ), .ip2(n19384), .s(
        n19368), .op(n9372) );
  mux2_1 U22203 ( .ip1(\pipeline/regfile/data[23][12] ), .ip2(n19384), .s(
        n19369), .op(n9180) );
  mux2_1 U22204 ( .ip1(\pipeline/regfile/data[12][12] ), .ip2(n19384), .s(
        n19370), .op(n9532) );
  mux2_1 U22205 ( .ip1(\pipeline/regfile/data[7][12] ), .ip2(n19384), .s(
        n19371), .op(n9692) );
  mux2_1 U22206 ( .ip1(\pipeline/regfile/data[8][12] ), .ip2(n19384), .s(
        n19372), .op(n9660) );
  mux2_1 U22207 ( .ip1(\pipeline/regfile/data[15][12] ), .ip2(n19384), .s(
        n19373), .op(n9436) );
  mux2_1 U22208 ( .ip1(\pipeline/regfile/data[10][12] ), .ip2(n19384), .s(
        n19374), .op(n9596) );
  mux2_1 U22209 ( .ip1(\pipeline/regfile/data[21][12] ), .ip2(n19384), .s(
        n19375), .op(n9244) );
  mux2_1 U22210 ( .ip1(\pipeline/regfile/data[24][12] ), .ip2(n19384), .s(
        n19376), .op(n9148) );
  mux2_1 U22211 ( .ip1(\pipeline/regfile/data[20][12] ), .ip2(n19384), .s(
        n19377), .op(n9276) );
  mux2_1 U22212 ( .ip1(\pipeline/regfile/data[9][12] ), .ip2(n19384), .s(
        n19378), .op(n9628) );
  mux2_1 U22213 ( .ip1(\pipeline/regfile/data[16][12] ), .ip2(n19384), .s(
        n19379), .op(n9404) );
  mux2_1 U22214 ( .ip1(\pipeline/regfile/data[3][12] ), .ip2(n19384), .s(
        n19380), .op(n9820) );
  mux2_1 U22215 ( .ip1(\pipeline/regfile/data[1][12] ), .ip2(n19384), .s(
        n19381), .op(n9884) );
  mux2_1 U22216 ( .ip1(\pipeline/regfile/data[2][12] ), .ip2(n19384), .s(
        n19382), .op(n9852) );
  mux2_1 U22217 ( .ip1(\pipeline/regfile/data[4][12] ), .ip2(n19384), .s(
        n19383), .op(n9788) );
  nand2_1 U22218 ( .ip1(n21238), .ip2(dmem_rdata[11]), .op(n19385) );
  or2_1 U22219 ( .ip1(n19385), .ip2(n22071), .op(n19389) );
  nand2_1 U22220 ( .ip1(n19386), .ip2(dmem_rdata[19]), .op(n19387) );
  or2_1 U22221 ( .ip1(n19387), .ip2(n22071), .op(n19388) );
  nand2_1 U22222 ( .ip1(n19389), .ip2(n19388), .op(n19391) );
  not_ab_or_c_or_d U22223 ( .ip1(n19392), .ip2(n21583), .ip3(n19391), .ip4(
        n19390), .op(n19394) );
  nand2_1 U22224 ( .ip1(dmem_rdata[27]), .ip2(n19410), .op(n19393) );
  nand2_1 U22225 ( .ip1(n19394), .ip2(n19393), .op(n19395) );
  mux2_1 U22226 ( .ip1(\pipeline/regfile/data[29][11] ), .ip2(n19395), .s(
        n21619), .op(n8989) );
  mux2_1 U22227 ( .ip1(\pipeline/regfile/data[14][11] ), .ip2(n19395), .s(
        n21604), .op(n9469) );
  mux2_1 U22228 ( .ip1(\pipeline/regfile/data[22][11] ), .ip2(n19395), .s(
        n21589), .op(n9213) );
  mux2_1 U22229 ( .ip1(\pipeline/regfile/data[5][11] ), .ip2(n19395), .s(
        n21598), .op(n9757) );
  mux2_1 U22230 ( .ip1(\pipeline/regfile/data[27][11] ), .ip2(n19395), .s(
        n21612), .op(n9053) );
  mux2_1 U22231 ( .ip1(\pipeline/regfile/data[26][11] ), .ip2(n19395), .s(
        n21607), .op(n9085) );
  mux2_1 U22232 ( .ip1(\pipeline/regfile/data[28][11] ), .ip2(n19395), .s(
        n21590), .op(n9021) );
  mux2_1 U22233 ( .ip1(\pipeline/regfile/data[31][11] ), .ip2(n19395), .s(
        n21606), .op(n8925) );
  mux2_1 U22234 ( .ip1(\pipeline/regfile/data[19][11] ), .ip2(n19395), .s(
        n21592), .op(n9309) );
  mux2_1 U22235 ( .ip1(\pipeline/regfile/data[6][11] ), .ip2(n19395), .s(
        n21597), .op(n9725) );
  mux2_1 U22236 ( .ip1(\pipeline/regfile/data[30][11] ), .ip2(n19395), .s(
        n21594), .op(n8957) );
  mux2_1 U22237 ( .ip1(\pipeline/regfile/data[18][11] ), .ip2(n19395), .s(
        n21595), .op(n9341) );
  mux2_1 U22238 ( .ip1(\pipeline/regfile/data[11][11] ), .ip2(n19395), .s(
        n21593), .op(n9565) );
  mux2_1 U22239 ( .ip1(\pipeline/regfile/data[25][11] ), .ip2(n19395), .s(
        n21602), .op(n9117) );
  mux2_1 U22240 ( .ip1(\pipeline/regfile/data[13][11] ), .ip2(n19395), .s(
        n21600), .op(n9501) );
  mux2_1 U22241 ( .ip1(\pipeline/regfile/data[17][11] ), .ip2(n19395), .s(
        n21616), .op(n9373) );
  mux2_1 U22242 ( .ip1(\pipeline/regfile/data[23][11] ), .ip2(n19395), .s(
        n21596), .op(n9181) );
  mux2_1 U22243 ( .ip1(\pipeline/regfile/data[12][11] ), .ip2(n19395), .s(
        n21591), .op(n9533) );
  mux2_1 U22244 ( .ip1(\pipeline/regfile/data[7][11] ), .ip2(n19395), .s(
        n21614), .op(n9693) );
  mux2_1 U22245 ( .ip1(\pipeline/regfile/data[8][11] ), .ip2(n19395), .s(
        n21617), .op(n9661) );
  mux2_1 U22246 ( .ip1(\pipeline/regfile/data[15][11] ), .ip2(n19395), .s(
        n21613), .op(n9437) );
  mux2_1 U22247 ( .ip1(\pipeline/regfile/data[10][11] ), .ip2(n19395), .s(
        n21618), .op(n9597) );
  mux2_1 U22248 ( .ip1(\pipeline/regfile/data[21][11] ), .ip2(n19395), .s(
        n21615), .op(n9245) );
  mux2_1 U22249 ( .ip1(\pipeline/regfile/data[24][11] ), .ip2(n19395), .s(
        n21603), .op(n9149) );
  mux2_1 U22250 ( .ip1(\pipeline/regfile/data[20][11] ), .ip2(n19395), .s(
        n21601), .op(n9277) );
  mux2_1 U22251 ( .ip1(\pipeline/regfile/data[9][11] ), .ip2(n19395), .s(
        n21609), .op(n9629) );
  mux2_1 U22252 ( .ip1(\pipeline/regfile/data[16][11] ), .ip2(n19395), .s(
        n21608), .op(n9405) );
  mux2_1 U22253 ( .ip1(\pipeline/regfile/data[3][11] ), .ip2(n19395), .s(
        n21599), .op(n9821) );
  mux2_1 U22254 ( .ip1(\pipeline/regfile/data[1][11] ), .ip2(n19395), .s(
        n21611), .op(n9885) );
  mux2_1 U22255 ( .ip1(\pipeline/regfile/data[2][11] ), .ip2(n19395), .s(
        n21610), .op(n9853) );
  mux2_1 U22256 ( .ip1(\pipeline/regfile/data[4][11] ), .ip2(n19395), .s(
        n21605), .op(n9789) );
  inv_1 U22257 ( .ip(n19396), .op(n19397) );
  nor2_1 U22258 ( .ip1(n19397), .ip2(n19404), .op(n19400) );
  nand2_1 U22259 ( .ip1(n21238), .ip2(dmem_rdata[10]), .op(n19398) );
  nor2_1 U22260 ( .ip1(n22071), .ip2(n19398), .op(n19399) );
  not_ab_or_c_or_d U22261 ( .ip1(n19409), .ip2(dmem_rdata[18]), .ip3(n19400), 
        .ip4(n19399), .op(n19402) );
  nand2_1 U22262 ( .ip1(n19410), .ip2(dmem_rdata[26]), .op(n19401) );
  nand3_1 U22263 ( .ip1(n19402), .ip2(n19412), .ip3(n19401), .op(n19403) );
  mux2_1 U22264 ( .ip1(\pipeline/regfile/data[29][10] ), .ip2(n19403), .s(
        n21619), .op(n8990) );
  mux2_1 U22265 ( .ip1(\pipeline/regfile/data[14][10] ), .ip2(n19403), .s(
        n21604), .op(n9470) );
  mux2_1 U22266 ( .ip1(\pipeline/regfile/data[22][10] ), .ip2(n19403), .s(
        n21589), .op(n9214) );
  mux2_1 U22267 ( .ip1(\pipeline/regfile/data[5][10] ), .ip2(n19403), .s(
        n21598), .op(n9758) );
  mux2_1 U22268 ( .ip1(\pipeline/regfile/data[27][10] ), .ip2(n19403), .s(
        n21612), .op(n9054) );
  mux2_1 U22269 ( .ip1(\pipeline/regfile/data[26][10] ), .ip2(n19403), .s(
        n21607), .op(n9086) );
  mux2_1 U22270 ( .ip1(\pipeline/regfile/data[28][10] ), .ip2(n19403), .s(
        n21590), .op(n9022) );
  mux2_1 U22271 ( .ip1(\pipeline/regfile/data[31][10] ), .ip2(n19403), .s(
        n21606), .op(n8926) );
  mux2_1 U22272 ( .ip1(\pipeline/regfile/data[19][10] ), .ip2(n19403), .s(
        n21592), .op(n9310) );
  mux2_1 U22273 ( .ip1(\pipeline/regfile/data[6][10] ), .ip2(n19403), .s(
        n21597), .op(n9726) );
  mux2_1 U22274 ( .ip1(\pipeline/regfile/data[30][10] ), .ip2(n19403), .s(
        n21594), .op(n8958) );
  mux2_1 U22275 ( .ip1(\pipeline/regfile/data[18][10] ), .ip2(n19403), .s(
        n21595), .op(n9342) );
  mux2_1 U22276 ( .ip1(\pipeline/regfile/data[11][10] ), .ip2(n19403), .s(
        n21593), .op(n9566) );
  mux2_1 U22277 ( .ip1(\pipeline/regfile/data[25][10] ), .ip2(n19403), .s(
        n21602), .op(n9118) );
  mux2_1 U22278 ( .ip1(\pipeline/regfile/data[13][10] ), .ip2(n19403), .s(
        n21600), .op(n9502) );
  mux2_1 U22279 ( .ip1(\pipeline/regfile/data[17][10] ), .ip2(n19403), .s(
        n21616), .op(n9374) );
  mux2_1 U22280 ( .ip1(\pipeline/regfile/data[23][10] ), .ip2(n19403), .s(
        n21596), .op(n9182) );
  mux2_1 U22281 ( .ip1(\pipeline/regfile/data[12][10] ), .ip2(n19403), .s(
        n21591), .op(n9534) );
  mux2_1 U22282 ( .ip1(\pipeline/regfile/data[7][10] ), .ip2(n19403), .s(
        n21614), .op(n9694) );
  mux2_1 U22283 ( .ip1(\pipeline/regfile/data[8][10] ), .ip2(n19403), .s(
        n21617), .op(n9662) );
  mux2_1 U22284 ( .ip1(\pipeline/regfile/data[15][10] ), .ip2(n19403), .s(
        n21613), .op(n9438) );
  mux2_1 U22285 ( .ip1(\pipeline/regfile/data[10][10] ), .ip2(n19403), .s(
        n21618), .op(n9598) );
  mux2_1 U22286 ( .ip1(\pipeline/regfile/data[21][10] ), .ip2(n19403), .s(
        n21615), .op(n9246) );
  mux2_1 U22287 ( .ip1(\pipeline/regfile/data[24][10] ), .ip2(n19403), .s(
        n21603), .op(n9150) );
  mux2_1 U22288 ( .ip1(\pipeline/regfile/data[20][10] ), .ip2(n19403), .s(
        n21601), .op(n9278) );
  mux2_1 U22289 ( .ip1(\pipeline/regfile/data[9][10] ), .ip2(n19403), .s(
        n21609), .op(n9630) );
  mux2_1 U22290 ( .ip1(\pipeline/regfile/data[16][10] ), .ip2(n19403), .s(
        n21608), .op(n9406) );
  mux2_1 U22291 ( .ip1(\pipeline/regfile/data[3][10] ), .ip2(n19403), .s(
        n21599), .op(n9822) );
  mux2_1 U22292 ( .ip1(\pipeline/regfile/data[1][10] ), .ip2(n19403), .s(
        n21611), .op(n9886) );
  mux2_1 U22293 ( .ip1(\pipeline/regfile/data[2][10] ), .ip2(n19403), .s(
        n21610), .op(n9854) );
  mux2_1 U22294 ( .ip1(\pipeline/regfile/data[4][10] ), .ip2(n19403), .s(
        n21605), .op(n9790) );
  nor2_1 U22295 ( .ip1(n19405), .ip2(n19404), .op(n19408) );
  nand2_1 U22296 ( .ip1(dmem_rdata[8]), .ip2(n21238), .op(n19406) );
  nor2_1 U22297 ( .ip1(n22071), .ip2(n19406), .op(n19407) );
  not_ab_or_c_or_d U22298 ( .ip1(n19409), .ip2(dmem_rdata[16]), .ip3(n19408), 
        .ip4(n19407), .op(n19413) );
  nand2_1 U22299 ( .ip1(n19410), .ip2(dmem_rdata[24]), .op(n19411) );
  nand3_1 U22300 ( .ip1(n19413), .ip2(n19412), .ip3(n19411), .op(n19414) );
  mux2_1 U22301 ( .ip1(\pipeline/regfile/data[29][8] ), .ip2(n19414), .s(
        n21619), .op(n8992) );
  mux2_1 U22302 ( .ip1(\pipeline/regfile/data[14][8] ), .ip2(n19414), .s(
        n21604), .op(n9472) );
  mux2_1 U22303 ( .ip1(\pipeline/regfile/data[22][8] ), .ip2(n19414), .s(
        n21589), .op(n9216) );
  mux2_1 U22304 ( .ip1(\pipeline/regfile/data[5][8] ), .ip2(n19414), .s(n21598), .op(n9760) );
  mux2_1 U22305 ( .ip1(\pipeline/regfile/data[27][8] ), .ip2(n19414), .s(
        n21612), .op(n9056) );
  mux2_1 U22306 ( .ip1(\pipeline/regfile/data[26][8] ), .ip2(n19414), .s(
        n21607), .op(n9088) );
  mux2_1 U22307 ( .ip1(\pipeline/regfile/data[28][8] ), .ip2(n19414), .s(
        n21590), .op(n9024) );
  mux2_1 U22308 ( .ip1(\pipeline/regfile/data[31][8] ), .ip2(n19414), .s(
        n21606), .op(n8928) );
  mux2_1 U22309 ( .ip1(\pipeline/regfile/data[19][8] ), .ip2(n19414), .s(
        n21592), .op(n9312) );
  mux2_1 U22310 ( .ip1(\pipeline/regfile/data[6][8] ), .ip2(n19414), .s(n21597), .op(n9728) );
  mux2_1 U22311 ( .ip1(\pipeline/regfile/data[30][8] ), .ip2(n19414), .s(
        n21594), .op(n8960) );
  mux2_1 U22312 ( .ip1(\pipeline/regfile/data[18][8] ), .ip2(n19414), .s(
        n21595), .op(n9344) );
  mux2_1 U22313 ( .ip1(\pipeline/regfile/data[11][8] ), .ip2(n19414), .s(
        n21593), .op(n9568) );
  mux2_1 U22314 ( .ip1(\pipeline/regfile/data[25][8] ), .ip2(n19414), .s(
        n21602), .op(n9120) );
  mux2_1 U22315 ( .ip1(\pipeline/regfile/data[13][8] ), .ip2(n19414), .s(
        n21600), .op(n9504) );
  mux2_1 U22316 ( .ip1(\pipeline/regfile/data[17][8] ), .ip2(n19414), .s(
        n21616), .op(n9376) );
  mux2_1 U22317 ( .ip1(\pipeline/regfile/data[23][8] ), .ip2(n19414), .s(
        n21596), .op(n9184) );
  mux2_1 U22318 ( .ip1(\pipeline/regfile/data[12][8] ), .ip2(n19414), .s(
        n21591), .op(n9536) );
  mux2_1 U22319 ( .ip1(\pipeline/regfile/data[7][8] ), .ip2(n19414), .s(n21614), .op(n9696) );
  mux2_1 U22320 ( .ip1(\pipeline/regfile/data[8][8] ), .ip2(n19414), .s(n21617), .op(n9664) );
  mux2_1 U22321 ( .ip1(\pipeline/regfile/data[15][8] ), .ip2(n19414), .s(
        n21613), .op(n9440) );
  mux2_1 U22322 ( .ip1(\pipeline/regfile/data[10][8] ), .ip2(n19414), .s(
        n21618), .op(n9600) );
  mux2_1 U22323 ( .ip1(\pipeline/regfile/data[21][8] ), .ip2(n19414), .s(
        n21615), .op(n9248) );
  mux2_1 U22324 ( .ip1(\pipeline/regfile/data[24][8] ), .ip2(n19414), .s(
        n21603), .op(n9152) );
  mux2_1 U22325 ( .ip1(\pipeline/regfile/data[20][8] ), .ip2(n19414), .s(
        n21601), .op(n9280) );
  mux2_1 U22326 ( .ip1(\pipeline/regfile/data[9][8] ), .ip2(n19414), .s(n21609), .op(n9632) );
  mux2_1 U22327 ( .ip1(\pipeline/regfile/data[16][8] ), .ip2(n19414), .s(
        n21608), .op(n9408) );
  mux2_1 U22328 ( .ip1(\pipeline/regfile/data[3][8] ), .ip2(n19414), .s(n21599), .op(n9824) );
  mux2_1 U22329 ( .ip1(\pipeline/regfile/data[1][8] ), .ip2(n19414), .s(n21611), .op(n9888) );
  mux2_1 U22330 ( .ip1(\pipeline/regfile/data[2][8] ), .ip2(n19414), .s(n21610), .op(n9856) );
  mux2_1 U22331 ( .ip1(\pipeline/regfile/data[4][8] ), .ip2(n19414), .s(n21605), .op(n9792) );
  nand2_1 U22332 ( .ip1(n19416), .ip2(n19415), .op(n19421) );
  nand2_1 U22333 ( .ip1(n20210), .ip2(n19417), .op(n19418) );
  nand2_1 U22334 ( .ip1(n19419), .ip2(n19418), .op(n19420) );
  xnor2_1 U22335 ( .ip1(n19421), .ip2(n19420), .op(n19448) );
  nor2_1 U22336 ( .ip1(n20887), .ip2(n19422), .op(n19425) );
  nor2_1 U22337 ( .ip1(n13881), .ip2(n19423), .op(n19424) );
  not_ab_or_c_or_d U22338 ( .ip1(n19427), .ip2(n19426), .ip3(n19425), .ip4(
        n19424), .op(n20882) );
  nor2_1 U22339 ( .ip1(n20724), .ip2(n20882), .op(n19447) );
  nand2_1 U22340 ( .ip1(n19428), .ip2(n21549), .op(n19445) );
  nand2_1 U22341 ( .ip1(n19429), .ip2(n19427), .op(n20227) );
  nor2_1 U22342 ( .ip1(n20894), .ip2(n20227), .op(n19437) );
  nand2_1 U22343 ( .ip1(n13636), .ip2(n19430), .op(n19431) );
  nand2_1 U22344 ( .ip1(n19431), .ip2(n21557), .op(n19435) );
  nand3_1 U22345 ( .ip1(n19433), .ip2(n20904), .ip3(n19432), .op(n19434) );
  nand3_1 U22346 ( .ip1(n19435), .ip2(n20735), .ip3(n19434), .op(n19436) );
  not_ab_or_c_or_d U22347 ( .ip1(n20911), .ip2(n19438), .ip3(n19437), .ip4(
        n19436), .op(n19444) );
  nand2_1 U22348 ( .ip1(n19440), .ip2(n19439), .op(n19443) );
  nand2_1 U22349 ( .ip1(n20231), .ip2(n19441), .op(n19442) );
  nand4_1 U22350 ( .ip1(n19445), .ip2(n19444), .ip3(n19443), .ip4(n19442), 
        .op(n19446) );
  ab_or_c_or_d U22351 ( .ip1(n19448), .ip2(n21577), .ip3(n19447), .ip4(n19446), 
        .op(dmem_haddr[15]) );
  mux2_1 U22352 ( .ip1(dmem_haddr[15]), .ip2(\pipeline/alu_out_WB [15]), .s(
        n21582), .op(n8717) );
  inv_1 U22353 ( .ip(n22177), .op(n19483) );
  nor2_1 U22354 ( .ip1(n19483), .ip2(n22267), .op(n19452) );
  not_ab_or_c_or_d U22355 ( .ip1(n19847), .ip2(n19450), .ip3(n19449), .ip4(
        n22276), .op(n19451) );
  or2_1 U22356 ( .ip1(n19452), .ip2(n19451), .op(\pipeline/csr/N1984 ) );
  inv_1 U22357 ( .ip(n19851), .op(n19453) );
  nor2_1 U22358 ( .ip1(\pipeline/csr/time_full [15]), .ip2(n19453), .op(n19455) );
  nor3_1 U22359 ( .ip1(n21177), .ip2(n19909), .ip3(n19455), .op(n19454) );
  not_ab_or_c_or_d U22360 ( .ip1(n21179), .ip2(n22177), .ip3(n21120), .ip4(
        n19454), .op(n19458) );
  nor2_1 U22361 ( .ip1(n19455), .ip2(n19909), .op(n19456) );
  nor2_1 U22362 ( .ip1(n22254), .ip2(n19456), .op(n19457) );
  nor2_1 U22363 ( .ip1(n19458), .ip2(n19457), .op(\pipeline/csr/N1952 ) );
  nand2_1 U22364 ( .ip1(n22008), .ip2(n22177), .op(n19461) );
  xor2_1 U22365 ( .ip1(n19860), .ip2(\pipeline/csr/mtime_full [15]), .op(
        n19459) );
  nand2_1 U22366 ( .ip1(n19459), .ip2(n22009), .op(n19460) );
  nand2_1 U22367 ( .ip1(n19461), .ip2(n19460), .op(\pipeline/csr/N2096 ) );
  nand2_1 U22368 ( .ip1(n22013), .ip2(\pipeline/csr/mscratch [15]), .op(n19463) );
  nand2_1 U22369 ( .ip1(n22014), .ip2(n22177), .op(n19462) );
  nand2_1 U22370 ( .ip1(n19463), .ip2(n19462), .op(n9913) );
  nand2_1 U22371 ( .ip1(n22372), .ip2(\pipeline/csr/from_host [15]), .op(
        n19465) );
  nand2_1 U22372 ( .ip1(n22373), .ip2(n22177), .op(n19464) );
  nand2_1 U22373 ( .ip1(n19465), .ip2(n19464), .op(n9945) );
  nand2_1 U22374 ( .ip1(n22378), .ip2(n22177), .op(n19467) );
  nand2_1 U22375 ( .ip1(n22376), .ip2(\pipeline/csr/to_host [15]), .op(n19466)
         );
  nand2_1 U22376 ( .ip1(n19467), .ip2(n19466), .op(n8757) );
  inv_1 U22377 ( .ip(n19872), .op(n19468) );
  nor2_1 U22378 ( .ip1(\pipeline/csr/cycle_full [15]), .ip2(n19468), .op(
        n19470) );
  nor3_1 U22379 ( .ip1(n19934), .ip2(n19470), .ip3(n21215), .op(n19469) );
  not_ab_or_c_or_d U22380 ( .ip1(n21076), .ip2(n22177), .ip3(n21120), .ip4(
        n19469), .op(n19473) );
  nor2_1 U22381 ( .ip1(n19470), .ip2(n19934), .op(n19471) );
  nor2_1 U22382 ( .ip1(n22254), .ip2(n19471), .op(n19472) );
  nor2_1 U22383 ( .ip1(n19473), .ip2(n19472), .op(\pipeline/csr/N1888 ) );
  nand2_1 U22384 ( .ip1(n22363), .ip2(\pipeline/csr/mtimecmp [15]), .op(n19475) );
  nand2_1 U22385 ( .ip1(n22365), .ip2(n22177), .op(n19474) );
  nand2_1 U22386 ( .ip1(n19475), .ip2(n19474), .op(n10007) );
  inv_1 U22387 ( .ip(\pipeline/csr/instret_full [15]), .op(n19478) );
  mux2_1 U22388 ( .ip1(n19478), .ip2(\pipeline/csr/instret_full [15]), .s(
        n19476), .op(n19477) );
  nor2_1 U22389 ( .ip1(n21005), .ip2(n19477), .op(n19480) );
  nor2_1 U22390 ( .ip1(n20990), .ip2(n19478), .op(n19479) );
  ab_or_c_or_d U22391 ( .ip1(n21019), .ip2(n22177), .ip3(n19480), .ip4(n19479), 
        .op(n10123) );
  nand2_1 U22392 ( .ip1(\pipeline/csr/mie [15]), .ip2(n22356), .op(n19482) );
  nand2_1 U22393 ( .ip1(n22357), .ip2(n22177), .op(n19481) );
  nand2_1 U22394 ( .ip1(n19482), .ip2(n19481), .op(n10045) );
  nor2_1 U22395 ( .ip1(n19483), .ip2(n22305), .op(n19486) );
  not_ab_or_c_or_d U22396 ( .ip1(n19889), .ip2(n19484), .ip3(n19952), .ip4(
        n22308), .op(n19485) );
  or2_1 U22397 ( .ip1(n19486), .ip2(n19485), .op(\pipeline/csr/N1920 ) );
  inv_1 U22398 ( .ip(n19487), .op(n19488) );
  mux2_1 U22399 ( .ip1(\pipeline/csr_rdata_WB [15]), .ip2(n19488), .s(n20389), 
        .op(n8791) );
  nor2_1 U22400 ( .ip1(n10183), .ip2(n20040), .op(n19493) );
  inv_1 U22401 ( .ip(n19490), .op(n20038) );
  xor2_1 U22402 ( .ip1(n19493), .ip2(n19492), .op(imem_haddr[20]) );
  nand2_1 U22403 ( .ip1(n21995), .ip2(imem_haddr[20]), .op(n19495) );
  nand2_1 U22404 ( .ip1(\pipeline/PC_IF [20]), .ip2(n21996), .op(n19494) );
  nand2_1 U22405 ( .ip1(n19495), .ip2(n19494), .op(n8450) );
  nand2_1 U22406 ( .ip1(\pipeline/PC_IF [20]), .ip2(n21988), .op(n19497) );
  nand2_1 U22407 ( .ip1(\pipeline/PC_DX [20]), .ip2(n21999), .op(n19496) );
  nand2_1 U22408 ( .ip1(n19497), .ip2(n19496), .op(n8449) );
  mux2_1 U22409 ( .ip1(\pipeline/PC_WB [20]), .ip2(\pipeline/PC_DX [20]), .s(
        n19498), .op(n8883) );
  nand2_1 U22410 ( .ip1(n19549), .ip2(n21043), .op(n19502) );
  xor2_1 U22411 ( .ip1(\pipeline/PC_WB [20]), .ip2(n20030), .op(n19499) );
  nand2_1 U22412 ( .ip1(n19499), .ip2(n21046), .op(n19501) );
  nand2_1 U22413 ( .ip1(n21174), .ip2(\pipeline/epc [20]), .op(n19500) );
  nand3_1 U22414 ( .ip1(n19502), .ip2(n19501), .ip3(n19500), .op(n8851) );
  nand2_1 U22415 ( .ip1(n21032), .ip2(n19549), .op(n19504) );
  nand2_1 U22416 ( .ip1(\pipeline/csr/mtvec [20]), .ip2(n20705), .op(n19503)
         );
  nand2_1 U22417 ( .ip1(n19504), .ip2(n19503), .op(n9972) );
  mux2_1 U22418 ( .ip1(dmem_haddr[20]), .ip2(\pipeline/alu_out_WB [20]), .s(
        n19505), .op(n8712) );
  inv_1 U22419 ( .ip(\pipeline/csr/time_full [52]), .op(n19507) );
  nor2_1 U22420 ( .ip1(n19508), .ip2(n19507), .op(n19506) );
  not_ab_or_c_or_d U22421 ( .ip1(n19508), .ip2(n19507), .ip3(n22282), .ip4(
        n19506), .op(n19511) );
  inv_1 U22422 ( .ip(n19549), .op(n22194) );
  nor2_1 U22423 ( .ip1(n22194), .ip2(n20748), .op(n19509) );
  nor2_1 U22424 ( .ip1(n19509), .ip2(n22284), .op(n19510) );
  nor2_1 U22425 ( .ip1(n19511), .ip2(n19510), .op(\pipeline/csr/N1989 ) );
  xnor2_1 U22426 ( .ip1(n19512), .ip2(\pipeline/csr/time_full [20]), .op(
        n19514) );
  nor2_1 U22427 ( .ip1(n21177), .ip2(n19514), .op(n19513) );
  not_ab_or_c_or_d U22428 ( .ip1(n21179), .ip2(n19549), .ip3(n21120), .ip4(
        n19513), .op(n19517) );
  inv_1 U22429 ( .ip(n19514), .op(n19515) );
  nor2_1 U22430 ( .ip1(n22254), .ip2(n19515), .op(n19516) );
  nor2_1 U22431 ( .ip1(n19517), .ip2(n19516), .op(\pipeline/csr/N1957 ) );
  inv_1 U22432 ( .ip(n19518), .op(n19519) );
  nor2_1 U22433 ( .ip1(\pipeline/csr/mtime_full [20]), .ip2(n19519), .op(
        n19522) );
  nor3_1 U22434 ( .ip1(n21193), .ip2(n19521), .ip3(n19522), .op(n19520) );
  not_ab_or_c_or_d U22435 ( .ip1(n21195), .ip2(n19549), .ip3(n21120), .ip4(
        n19520), .op(n19525) );
  nor2_1 U22436 ( .ip1(n19522), .ip2(n19521), .op(n19523) );
  nor2_1 U22437 ( .ip1(n22254), .ip2(n19523), .op(n19524) );
  nor2_1 U22438 ( .ip1(n19525), .ip2(n19524), .op(\pipeline/csr/N2101 ) );
  nand2_1 U22439 ( .ip1(\pipeline/csr/mscratch [20]), .ip2(n22013), .op(n19527) );
  nand2_1 U22440 ( .ip1(n22014), .ip2(n19549), .op(n19526) );
  nand2_1 U22441 ( .ip1(n19527), .ip2(n19526), .op(n9908) );
  nand2_1 U22442 ( .ip1(\pipeline/csr/from_host [20]), .ip2(n22372), .op(
        n19529) );
  nand2_1 U22443 ( .ip1(n22373), .ip2(n19549), .op(n19528) );
  nand2_1 U22444 ( .ip1(n19529), .ip2(n19528), .op(n9940) );
  nand2_1 U22445 ( .ip1(n22378), .ip2(n19549), .op(n19531) );
  nand2_1 U22446 ( .ip1(\pipeline/csr/to_host [20]), .ip2(n22376), .op(n19530)
         );
  nand2_1 U22447 ( .ip1(n19531), .ip2(n19530), .op(n8752) );
  or2_1 U22448 ( .ip1(\pipeline/csr/cycle_full [20]), .ip2(n19532), .op(n19533) );
  nand2_1 U22449 ( .ip1(n19534), .ip2(n19533), .op(n19535) );
  or2_1 U22450 ( .ip1(n21145), .ip2(n19535), .op(n19537) );
  nand2_1 U22451 ( .ip1(n22021), .ip2(n19549), .op(n19536) );
  nand2_1 U22452 ( .ip1(n19537), .ip2(n19536), .op(\pipeline/csr/N1893 ) );
  nand2_1 U22453 ( .ip1(\pipeline/csr/mtimecmp [20]), .ip2(n22363), .op(n19539) );
  nand2_1 U22454 ( .ip1(n22365), .ip2(n19549), .op(n19538) );
  nand2_1 U22455 ( .ip1(n19539), .ip2(n19538), .op(n10002) );
  nand2_1 U22456 ( .ip1(n21019), .ip2(n19549), .op(n19546) );
  nand2_1 U22457 ( .ip1(\pipeline/csr/instret_full [20]), .ip2(n21016), .op(
        n19545) );
  mux2_1 U22458 ( .ip1(\pipeline/csr/instret_full [20]), .ip2(n19541), .s(
        n19540), .op(n19543) );
  nor2_1 U22459 ( .ip1(n21012), .ip2(n21011), .op(n19542) );
  or2_1 U22460 ( .ip1(n19543), .ip2(n19542), .op(n19544) );
  nand3_1 U22461 ( .ip1(n19546), .ip2(n19545), .ip3(n19544), .op(n10118) );
  nand2_1 U22462 ( .ip1(\pipeline/csr/mie [20]), .ip2(n22356), .op(n19548) );
  nand2_1 U22463 ( .ip1(n22357), .ip2(n19549), .op(n19547) );
  nand2_1 U22464 ( .ip1(n19548), .ip2(n19547), .op(n10040) );
  nand2_1 U22465 ( .ip1(n22314), .ip2(n19549), .op(n19554) );
  or2_1 U22466 ( .ip1(\pipeline/csr/cycle_full [52]), .ip2(n19550), .op(n19551) );
  nand3_1 U22467 ( .ip1(n19552), .ip2(n19551), .ip3(n22316), .op(n19553) );
  nand2_1 U22468 ( .ip1(n19554), .ip2(n19553), .op(\pipeline/csr/N1925 ) );
  inv_1 U22469 ( .ip(n19555), .op(n19556) );
  mux2_1 U22470 ( .ip1(\pipeline/csr_rdata_WB [20]), .ip2(n19556), .s(n22067), 
        .op(n8786) );
  nand2_1 U22471 ( .ip1(imem_haddr[24]), .ip2(n21995), .op(n19558) );
  nand2_1 U22472 ( .ip1(\pipeline/PC_IF [24]), .ip2(n21996), .op(n19557) );
  nand2_1 U22473 ( .ip1(n19558), .ip2(n19557), .op(n8442) );
  nand2_1 U22474 ( .ip1(\pipeline/PC_IF [24]), .ip2(n22048), .op(n19560) );
  nand2_1 U22475 ( .ip1(\pipeline/PC_DX [24]), .ip2(n21999), .op(n19559) );
  nand2_1 U22476 ( .ip1(n19560), .ip2(n19559), .op(n8441) );
  mux2_1 U22477 ( .ip1(dmem_haddr[7]), .ip2(\pipeline/alu_out_WB [7]), .s(
        n21582), .op(n8725) );
  inv_1 U22478 ( .ip(n19677), .op(n19680) );
  nor2_1 U22479 ( .ip1(n19680), .ip2(n22267), .op(n19563) );
  not_ab_or_c_or_d U22480 ( .ip1(n20330), .ip2(n19561), .ip3(n19695), .ip4(
        n22276), .op(n19562) );
  or2_1 U22481 ( .ip1(n19563), .ip2(n19562), .op(\pipeline/csr/N1976 ) );
  inv_1 U22482 ( .ip(n20344), .op(n19564) );
  nor2_1 U22483 ( .ip1(\pipeline/csr/time_full [7]), .ip2(n19564), .op(n19566)
         );
  nor3_1 U22484 ( .ip1(n21177), .ip2(n19702), .ip3(n19566), .op(n19565) );
  not_ab_or_c_or_d U22485 ( .ip1(n21179), .ip2(n19677), .ip3(n21217), .ip4(
        n19565), .op(n19569) );
  nor2_1 U22486 ( .ip1(n19566), .ip2(n19702), .op(n19567) );
  nor2_1 U22487 ( .ip1(n22254), .ip2(n19567), .op(n19568) );
  nor2_1 U22488 ( .ip1(n19569), .ip2(n19568), .op(\pipeline/csr/N1944 ) );
  nand2_1 U22489 ( .ip1(n22008), .ip2(n19677), .op(n19572) );
  xor2_1 U22490 ( .ip1(\pipeline/csr/mtime_full [7]), .ip2(n20353), .op(n19570) );
  nand2_1 U22491 ( .ip1(n19570), .ip2(n22009), .op(n19571) );
  nand2_1 U22492 ( .ip1(n19572), .ip2(n19571), .op(\pipeline/csr/N2088 ) );
  nand2_1 U22493 ( .ip1(\pipeline/csr/mscratch [7]), .ip2(n22013), .op(n19574)
         );
  nand2_1 U22494 ( .ip1(n22014), .ip2(n19677), .op(n19573) );
  nand2_1 U22495 ( .ip1(n19574), .ip2(n19573), .op(n9921) );
  nand2_1 U22496 ( .ip1(\pipeline/csr/from_host [7]), .ip2(n22372), .op(n19576) );
  nand2_1 U22497 ( .ip1(n22373), .ip2(n19677), .op(n19575) );
  nand2_1 U22498 ( .ip1(n19576), .ip2(n19575), .op(n9953) );
  nand2_1 U22499 ( .ip1(n22378), .ip2(n19677), .op(n19578) );
  nand2_1 U22500 ( .ip1(\pipeline/csr/to_host [7]), .ip2(n22376), .op(n19577)
         );
  nand2_1 U22501 ( .ip1(n19578), .ip2(n19577), .op(n8765) );
  xor2_1 U22502 ( .ip1(\pipeline/csr/mtime_full [39]), .ip2(n22151), .op(
        n19579) );
  nand2_1 U22503 ( .ip1(n19579), .ip2(n18449), .op(n19581) );
  nand2_1 U22504 ( .ip1(n22235), .ip2(n19677), .op(n19580) );
  nand2_1 U22505 ( .ip1(n19581), .ip2(n19580), .op(\pipeline/csr/N2120 ) );
  inv_1 U22506 ( .ip(n20365), .op(n19582) );
  nor2_1 U22507 ( .ip1(\pipeline/csr/cycle_full [7]), .ip2(n19582), .op(n19584) );
  nor3_1 U22508 ( .ip1(n19729), .ip2(n19584), .ip3(n21215), .op(n19583) );
  not_ab_or_c_or_d U22509 ( .ip1(n21076), .ip2(n19677), .ip3(n21120), .ip4(
        n19583), .op(n19587) );
  nor2_1 U22510 ( .ip1(n19584), .ip2(n19729), .op(n19585) );
  nor2_1 U22511 ( .ip1(n22254), .ip2(n19585), .op(n19586) );
  nor2_1 U22512 ( .ip1(n19587), .ip2(n19586), .op(\pipeline/csr/N1880 ) );
  nand2_1 U22513 ( .ip1(\pipeline/csr/mtimecmp [7]), .ip2(n22363), .op(n19589)
         );
  nand2_1 U22514 ( .ip1(n22365), .ip2(n19677), .op(n19588) );
  nand2_1 U22515 ( .ip1(n19589), .ip2(n19588), .op(n10015) );
  nor2_1 U22516 ( .ip1(n19680), .ip2(n21001), .op(n19593) );
  inv_1 U22517 ( .ip(\pipeline/csr/instret_full [7]), .op(n19590) );
  mux2_1 U22518 ( .ip1(n19590), .ip2(\pipeline/csr/instret_full [7]), .s(
        n20369), .op(n19591) );
  nor2_1 U22519 ( .ip1(n21005), .ip2(n19591), .op(n19592) );
  ab_or_c_or_d U22520 ( .ip1(n21016), .ip2(\pipeline/csr/instret_full [7]), 
        .ip3(n19593), .ip4(n19592), .op(n10131) );
  nand2_1 U22521 ( .ip1(\pipeline/csr/mie [7]), .ip2(n22356), .op(n19595) );
  nand2_1 U22522 ( .ip1(n22357), .ip2(n19677), .op(n19594) );
  nand2_1 U22523 ( .ip1(n19595), .ip2(n19594), .op(n10053) );
  nor2_1 U22524 ( .ip1(n19680), .ip2(n22305), .op(n19598) );
  not_ab_or_c_or_d U22525 ( .ip1(n20375), .ip2(n19596), .ip3(n19740), .ip4(
        n22308), .op(n19597) );
  or2_1 U22526 ( .ip1(n19598), .ip2(n19597), .op(\pipeline/csr/N1912 ) );
  inv_1 U22527 ( .ip(n19599), .op(n19600) );
  nor2_1 U22528 ( .ip1(n19601), .ip2(n19600), .op(n21231) );
  inv_1 U22529 ( .ip(n21231), .op(n19676) );
  inv_1 U22530 ( .ip(\pipeline/csr/mtime_full [19]), .op(n19602) );
  mux2_1 U22531 ( .ip1(n19602), .ip2(\pipeline/csr/mtime_full [19]), .s(
        \pipeline/csr/mtimecmp [19]), .op(n19609) );
  inv_1 U22532 ( .ip(\pipeline/csr/mtime_full [9]), .op(n19603) );
  mux2_1 U22533 ( .ip1(n19603), .ip2(\pipeline/csr/mtime_full [9]), .s(
        \pipeline/csr/mtimecmp [9]), .op(n19608) );
  mux2_1 U22534 ( .ip1(n19604), .ip2(\pipeline/csr/mtime_full [22]), .s(
        \pipeline/csr/mtimecmp [22]), .op(n19607) );
  inv_1 U22535 ( .ip(\pipeline/csr/mtime_full [13]), .op(n19605) );
  mux2_1 U22536 ( .ip1(n19605), .ip2(\pipeline/csr/mtime_full [13]), .s(
        \pipeline/csr/mtimecmp [13]), .op(n19606) );
  nand4_1 U22537 ( .ip1(n19609), .ip2(n19608), .ip3(n19607), .ip4(n19606), 
        .op(n19673) );
  mux2_1 U22538 ( .ip1(n19610), .ip2(\pipeline/csr/mtime_full [18]), .s(
        \pipeline/csr/mtimecmp [18]), .op(n19617) );
  mux2_1 U22539 ( .ip1(n19611), .ip2(\pipeline/csr/mtime_full [15]), .s(
        \pipeline/csr/mtimecmp [15]), .op(n19616) );
  inv_1 U22540 ( .ip(\pipeline/csr/mtime_full [7]), .op(n19612) );
  mux2_1 U22541 ( .ip1(n19612), .ip2(\pipeline/csr/mtime_full [7]), .s(
        \pipeline/csr/mtimecmp [7]), .op(n19615) );
  mux2_1 U22542 ( .ip1(n19613), .ip2(\pipeline/csr/mtime_full [27]), .s(
        \pipeline/csr/mtimecmp [27]), .op(n19614) );
  nand4_1 U22543 ( .ip1(n19617), .ip2(n19616), .ip3(n19615), .ip4(n19614), 
        .op(n19672) );
  mux2_1 U22544 ( .ip1(\pipeline/csr/mtime_full [3]), .ip2(n21191), .s(
        \pipeline/csr/mtimecmp [3]), .op(n19619) );
  nor2_1 U22545 ( .ip1(\pipeline/csr/mtimecmp [28]), .ip2(n19620), .op(n19618)
         );
  not_ab_or_c_or_d U22546 ( .ip1(\pipeline/csr/mtimecmp [28]), .ip2(n19620), 
        .ip3(n19619), .ip4(n19618), .op(n19634) );
  mux2_1 U22547 ( .ip1(\pipeline/csr/mtime_full [24]), .ip2(n19621), .s(
        \pipeline/csr/mtimecmp [24]), .op(n19628) );
  mux2_1 U22548 ( .ip1(\pipeline/csr/mtime_full [4]), .ip2(n19622), .s(
        \pipeline/csr/mtimecmp [4]), .op(n19627) );
  mux2_1 U22549 ( .ip1(\pipeline/csr/mtime_full [2]), .ip2(n19623), .s(
        \pipeline/csr/mtimecmp [2]), .op(n19626) );
  inv_1 U22550 ( .ip(\pipeline/csr/mtime_full [31]), .op(n19624) );
  mux2_1 U22551 ( .ip1(\pipeline/csr/mtime_full [31]), .ip2(n19624), .s(
        \pipeline/csr/mtimecmp [31]), .op(n19625) );
  nor4_1 U22552 ( .ip1(n19628), .ip2(n19627), .ip3(n19626), .ip4(n19625), .op(
        n19633) );
  mux2_1 U22553 ( .ip1(n19629), .ip2(\pipeline/csr/mtime_full [16]), .s(
        \pipeline/csr/mtimecmp [16]), .op(n19632) );
  mux2_1 U22554 ( .ip1(n19630), .ip2(\pipeline/csr/mtime_full [12]), .s(
        \pipeline/csr/mtimecmp [12]), .op(n19631) );
  nand4_1 U22555 ( .ip1(n19634), .ip2(n19633), .ip3(n19632), .ip4(n19631), 
        .op(n19671) );
  mux2_1 U22556 ( .ip1(\pipeline/csr/mtime_full [1]), .ip2(n19635), .s(
        \pipeline/csr/mtimecmp [1]), .op(n19642) );
  mux2_1 U22557 ( .ip1(\pipeline/csr/mtime_full [10]), .ip2(n19636), .s(
        \pipeline/csr/mtimecmp [10]), .op(n19641) );
  mux2_1 U22558 ( .ip1(\pipeline/csr/mtime_full [8]), .ip2(n19637), .s(
        \pipeline/csr/mtimecmp [8]), .op(n19640) );
  mux2_1 U22559 ( .ip1(\pipeline/csr/mtime_full [30]), .ip2(n19638), .s(
        \pipeline/csr/mtimecmp [30]), .op(n19639) );
  nor4_1 U22560 ( .ip1(n19642), .ip2(n19641), .ip3(n19640), .ip4(n19639), .op(
        n19669) );
  inv_1 U22561 ( .ip(\pipeline/csr/mtime_full [5]), .op(n19643) );
  mux2_1 U22562 ( .ip1(\pipeline/csr/mtime_full [5]), .ip2(n19643), .s(
        \pipeline/csr/mtimecmp [5]), .op(n19649) );
  inv_1 U22563 ( .ip(\pipeline/csr/mtime_full [23]), .op(n19644) );
  mux2_1 U22564 ( .ip1(\pipeline/csr/mtime_full [23]), .ip2(n19644), .s(
        \pipeline/csr/mtimecmp [23]), .op(n19648) );
  mux2_1 U22565 ( .ip1(\pipeline/csr/mtime_full [0]), .ip2(n20980), .s(
        \pipeline/csr/mtimecmp [0]), .op(n19647) );
  inv_1 U22566 ( .ip(\pipeline/csr/mtime_full [17]), .op(n19645) );
  mux2_1 U22567 ( .ip1(\pipeline/csr/mtime_full [17]), .ip2(n19645), .s(
        \pipeline/csr/mtimecmp [17]), .op(n19646) );
  nor4_1 U22568 ( .ip1(n19649), .ip2(n19648), .ip3(n19647), .ip4(n19646), .op(
        n19668) );
  mux2_1 U22569 ( .ip1(\pipeline/csr/mtime_full [14]), .ip2(n19650), .s(
        \pipeline/csr/mtimecmp [14]), .op(n19657) );
  inv_1 U22570 ( .ip(\pipeline/csr/mtime_full [11]), .op(n19651) );
  mux2_1 U22571 ( .ip1(\pipeline/csr/mtime_full [11]), .ip2(n19651), .s(
        \pipeline/csr/mtimecmp [11]), .op(n19656) );
  inv_1 U22572 ( .ip(\pipeline/csr/mtime_full [29]), .op(n19652) );
  mux2_1 U22573 ( .ip1(\pipeline/csr/mtime_full [29]), .ip2(n19652), .s(
        \pipeline/csr/mtimecmp [29]), .op(n19655) );
  inv_1 U22574 ( .ip(\pipeline/csr/mtime_full [25]), .op(n19653) );
  mux2_1 U22575 ( .ip1(\pipeline/csr/mtime_full [25]), .ip2(n19653), .s(
        \pipeline/csr/mtimecmp [25]), .op(n19654) );
  nor4_1 U22576 ( .ip1(n19657), .ip2(n19656), .ip3(n19655), .ip4(n19654), .op(
        n19667) );
  mux2_1 U22577 ( .ip1(\pipeline/csr/mtime_full [20]), .ip2(n19658), .s(
        \pipeline/csr/mtimecmp [20]), .op(n19665) );
  mux2_1 U22578 ( .ip1(\pipeline/csr/mtime_full [6]), .ip2(n19659), .s(
        \pipeline/csr/mtimecmp [6]), .op(n19664) );
  mux2_1 U22579 ( .ip1(\pipeline/csr/mtime_full [26]), .ip2(n19660), .s(
        \pipeline/csr/mtimecmp [26]), .op(n19663) );
  mux2_1 U22580 ( .ip1(\pipeline/csr/mtime_full [21]), .ip2(n19661), .s(
        \pipeline/csr/mtimecmp [21]), .op(n19662) );
  nor4_1 U22581 ( .ip1(n19665), .ip2(n19664), .ip3(n19663), .ip4(n19662), .op(
        n19666) );
  nand4_1 U22582 ( .ip1(n19669), .ip2(n19668), .ip3(n19667), .ip4(n19666), 
        .op(n19670) );
  nor4_1 U22583 ( .ip1(n19673), .ip2(n19672), .ip3(n19671), .ip4(n19670), .op(
        n19674) );
  or2_1 U22584 ( .ip1(\pipeline/csr/mip[7] ), .ip2(n19674), .op(n19675) );
  nand3_1 U22585 ( .ip1(n22363), .ip2(n19676), .ip3(n19675), .op(n19679) );
  nand3_1 U22586 ( .ip1(n21231), .ip2(n20966), .ip3(n19677), .op(n19678) );
  nand2_1 U22587 ( .ip1(n19679), .ip2(n19678), .op(n10073) );
  nor2_1 U22588 ( .ip1(n19680), .ip2(n21168), .op(n19686) );
  inv_1 U22589 ( .ip(\pipeline/PC_WB [7]), .op(n19684) );
  nand2_1 U22590 ( .ip1(n19681), .ip2(\pipeline/PC_WB [6]), .op(n19683) );
  not_ab_or_c_or_d U22591 ( .ip1(n19684), .ip2(n19683), .ip3(n19682), .ip4(
        n21171), .op(n19685) );
  ab_or_c_or_d U22592 ( .ip1(n21174), .ip2(\pipeline/epc [7]), .ip3(n19686), 
        .ip4(n19685), .op(n8864) );
  nor2_1 U22593 ( .ip1(n19688), .ip2(n14269), .op(n19690) );
  xor2_1 U22594 ( .ip1(n19690), .ip2(n19689), .op(imem_haddr[8]) );
  nand2_1 U22595 ( .ip1(n21995), .ip2(imem_haddr[8]), .op(n19692) );
  nand2_1 U22596 ( .ip1(\pipeline/PC_IF [8]), .ip2(n21996), .op(n19691) );
  nand2_1 U22597 ( .ip1(n19692), .ip2(n19691), .op(n8474) );
  nand2_1 U22598 ( .ip1(\pipeline/PC_IF [8]), .ip2(n21988), .op(n19694) );
  nand2_1 U22599 ( .ip1(\pipeline/PC_DX [8]), .ip2(n21999), .op(n19693) );
  nand2_1 U22600 ( .ip1(n19694), .ip2(n19693), .op(n8473) );
  mux2_1 U22601 ( .ip1(\pipeline/PC_WB [8]), .ip2(\pipeline/PC_DX [8]), .s(
        n17777), .op(n8895) );
  mux2_1 U22602 ( .ip1(dmem_haddr[8]), .ip2(\pipeline/alu_out_WB [8]), .s(
        n21582), .op(n8724) );
  nand2_1 U22603 ( .ip1(n22282), .ip2(n19739), .op(n19699) );
  or2_1 U22604 ( .ip1(\pipeline/csr/time_full [40]), .ip2(n19695), .op(n19696)
         );
  nand3_1 U22605 ( .ip1(n19697), .ip2(n19696), .ip3(n22284), .op(n19698) );
  nand2_1 U22606 ( .ip1(n19699), .ip2(n19698), .op(\pipeline/csr/N1977 ) );
  nand2_1 U22607 ( .ip1(n19700), .ip2(n22257), .op(n19701) );
  nand2_1 U22608 ( .ip1(n20181), .ip2(n19701), .op(n19705) );
  nand2_1 U22609 ( .ip1(n19705), .ip2(n21177), .op(n19704) );
  xor2_1 U22610 ( .ip1(\pipeline/csr/time_full [8]), .ip2(n19702), .op(n19703)
         );
  nand2_1 U22611 ( .ip1(n19704), .ip2(n19703), .op(n19707) );
  or2_1 U22612 ( .ip1(n21210), .ip2(n19705), .op(n19706) );
  nand2_1 U22613 ( .ip1(n19707), .ip2(n19706), .op(\pipeline/csr/N1945 ) );
  inv_1 U22614 ( .ip(n19708), .op(n19709) );
  nor2_1 U22615 ( .ip1(\pipeline/csr/mtime_full [8]), .ip2(n19709), .op(n19712) );
  nor3_1 U22616 ( .ip1(n21193), .ip2(n19712), .ip3(n19711), .op(n19710) );
  not_ab_or_c_or_d U22617 ( .ip1(n21195), .ip2(n19739), .ip3(n21120), .ip4(
        n19710), .op(n19715) );
  nor2_1 U22618 ( .ip1(n19712), .ip2(n19711), .op(n19713) );
  nor2_1 U22619 ( .ip1(n22254), .ip2(n19713), .op(n19714) );
  nor2_1 U22620 ( .ip1(n19715), .ip2(n19714), .op(\pipeline/csr/N2089 ) );
  nand2_1 U22621 ( .ip1(\pipeline/csr/mscratch [8]), .ip2(n22013), .op(n19717)
         );
  nand2_1 U22622 ( .ip1(n22014), .ip2(n19739), .op(n19716) );
  nand2_1 U22623 ( .ip1(n19717), .ip2(n19716), .op(n9920) );
  nand2_1 U22624 ( .ip1(\pipeline/csr/from_host [8]), .ip2(n22372), .op(n19719) );
  nand2_1 U22625 ( .ip1(n22373), .ip2(n19739), .op(n19718) );
  nand2_1 U22626 ( .ip1(n19719), .ip2(n19718), .op(n9952) );
  nand2_1 U22627 ( .ip1(n22378), .ip2(n19739), .op(n19721) );
  nand2_1 U22628 ( .ip1(\pipeline/csr/to_host [8]), .ip2(n22376), .op(n19720)
         );
  nand2_1 U22629 ( .ip1(n19721), .ip2(n19720), .op(n8764) );
  nand2_1 U22630 ( .ip1(n22235), .ip2(n19739), .op(n19728) );
  nor2_1 U22631 ( .ip1(n22247), .ip2(n19722), .op(n19726) );
  inv_1 U22632 ( .ip(n19723), .op(n19724) );
  or2_1 U22633 ( .ip1(\pipeline/csr/mtime_full [40]), .ip2(n19724), .op(n19725) );
  nand2_1 U22634 ( .ip1(n19726), .ip2(n19725), .op(n19727) );
  nand2_1 U22635 ( .ip1(n19728), .ip2(n19727), .op(\pipeline/csr/N2121 ) );
  or2_1 U22636 ( .ip1(\pipeline/csr/cycle_full [8]), .ip2(n19729), .op(n19730)
         );
  nand2_1 U22637 ( .ip1(n19731), .ip2(n19730), .op(n19732) );
  or2_1 U22638 ( .ip1(n21145), .ip2(n19732), .op(n19734) );
  nand2_1 U22639 ( .ip1(n22021), .ip2(n19739), .op(n19733) );
  nand2_1 U22640 ( .ip1(n19734), .ip2(n19733), .op(\pipeline/csr/N1881 ) );
  nand2_1 U22641 ( .ip1(\pipeline/csr/mtimecmp [8]), .ip2(n22363), .op(n19736)
         );
  nand2_1 U22642 ( .ip1(n22365), .ip2(n19739), .op(n19735) );
  nand2_1 U22643 ( .ip1(n19736), .ip2(n19735), .op(n10014) );
  nand2_1 U22644 ( .ip1(\pipeline/csr/mie [8]), .ip2(n22356), .op(n19738) );
  nand2_1 U22645 ( .ip1(n22357), .ip2(n19739), .op(n19737) );
  nand2_1 U22646 ( .ip1(n19738), .ip2(n19737), .op(n10052) );
  nand2_1 U22647 ( .ip1(n22314), .ip2(n19739), .op(n19744) );
  or2_1 U22648 ( .ip1(\pipeline/csr/cycle_full [40]), .ip2(n19740), .op(n19741) );
  nand3_1 U22649 ( .ip1(n19742), .ip2(n19741), .ip3(n22316), .op(n19743) );
  nand2_1 U22650 ( .ip1(n19744), .ip2(n19743), .op(\pipeline/csr/N1913 ) );
  inv_1 U22651 ( .ip(n19745), .op(n19746) );
  mux2_1 U22652 ( .ip1(\pipeline/csr_rdata_WB [8]), .ip2(n19746), .s(n17429), 
        .op(n8798) );
  xor2_1 U22653 ( .ip1(n19748), .ip2(n19747), .op(n19749) );
  nand2_1 U22654 ( .ip1(n21649), .ip2(n19749), .op(n19761) );
  inv_1 U22655 ( .ip(n19750), .op(n19751) );
  nand2_1 U22656 ( .ip1(n19752), .ip2(n19751), .op(n20384) );
  nand2_1 U22657 ( .ip1(n20384), .ip2(n19753), .op(n19754) );
  nand2_1 U22658 ( .ip1(n19755), .ip2(n19754), .op(n20496) );
  xor2_1 U22659 ( .ip1(n20496), .ip2(n19756), .op(n19757) );
  nor2_1 U22660 ( .ip1(n21884), .ip2(n19757), .op(n19758) );
  xor2_1 U22661 ( .ip1(\pipeline/md/a [8]), .ip2(n19758), .op(n19759) );
  nand2_1 U22662 ( .ip1(n19759), .ip2(n21643), .op(n19760) );
  nand2_1 U22663 ( .ip1(n19761), .ip2(n19760), .op(n8407) );
  mux2_1 U22664 ( .ip1(\pipeline/csr_rdata_WB [9]), .ip2(n19762), .s(n17777), 
        .op(n8797) );
  xor2_1 U22665 ( .ip1(n19764), .ip2(n19763), .op(imem_haddr[9]) );
  nor2_1 U22666 ( .ip1(\pipeline/PC_IF [9]), .ip2(n19765), .op(n19768) );
  nor2_1 U22667 ( .ip1(imem_haddr[9]), .ip2(n19766), .op(n19767) );
  nor2_1 U22668 ( .ip1(n19768), .ip2(n19767), .op(n8472) );
  nand2_1 U22669 ( .ip1(\pipeline/PC_IF [9]), .ip2(n21988), .op(n19770) );
  nand2_1 U22670 ( .ip1(\pipeline/PC_DX [9]), .ip2(n21999), .op(n19769) );
  nand2_1 U22671 ( .ip1(n19770), .ip2(n19769), .op(n8471) );
  mux2_1 U22672 ( .ip1(\pipeline/PC_WB [9]), .ip2(\pipeline/PC_DX [9]), .s(
        n19498), .op(n8894) );
  mux2_1 U22673 ( .ip1(\pipeline/PC_WB [10]), .ip2(\pipeline/PC_DX [10]), .s(
        n17777), .op(n8893) );
  nor2_1 U22674 ( .ip1(n19805), .ip2(n21168), .op(n19777) );
  inv_1 U22675 ( .ip(\pipeline/PC_WB [10]), .op(n19775) );
  inv_1 U22676 ( .ip(n19771), .op(n19772) );
  nand2_1 U22677 ( .ip1(n19772), .ip2(\pipeline/PC_WB [9]), .op(n19774) );
  not_ab_or_c_or_d U22678 ( .ip1(n19775), .ip2(n19774), .ip3(n19773), .ip4(
        n21171), .op(n19776) );
  ab_or_c_or_d U22679 ( .ip1(n21174), .ip2(\pipeline/epc [10]), .ip3(n19777), 
        .ip4(n19776), .op(n8861) );
  nand2_1 U22680 ( .ip1(n21032), .ip2(n19828), .op(n19779) );
  nand2_1 U22681 ( .ip1(\pipeline/csr/mtvec [10]), .ip2(n20705), .op(n19778)
         );
  nand2_1 U22682 ( .ip1(n19779), .ip2(n19778), .op(n9982) );
  mux2_1 U22683 ( .ip1(dmem_haddr[10]), .ip2(\pipeline/alu_out_WB [10]), .s(
        n19505), .op(n8722) );
  nand2_1 U22684 ( .ip1(n22282), .ip2(n19828), .op(n19783) );
  or2_1 U22685 ( .ip1(\pipeline/csr/time_full [42]), .ip2(n19780), .op(n19781)
         );
  nand3_1 U22686 ( .ip1(n20175), .ip2(n19781), .ip3(n22284), .op(n19782) );
  nand2_1 U22687 ( .ip1(n19783), .ip2(n19782), .op(\pipeline/csr/N1979 ) );
  or2_1 U22688 ( .ip1(\pipeline/csr/time_full [10]), .ip2(n19784), .op(n19785)
         );
  nand2_1 U22689 ( .ip1(n20183), .ip2(n19785), .op(n19787) );
  nor2_1 U22690 ( .ip1(n21177), .ip2(n19787), .op(n19786) );
  not_ab_or_c_or_d U22691 ( .ip1(n21179), .ip2(n19828), .ip3(n21120), .ip4(
        n19786), .op(n19790) );
  inv_1 U22692 ( .ip(n19787), .op(n19788) );
  nor2_1 U22693 ( .ip1(n22254), .ip2(n19788), .op(n19789) );
  nor2_1 U22694 ( .ip1(n19790), .ip2(n19789), .op(\pipeline/csr/N1947 ) );
  inv_1 U22695 ( .ip(n19791), .op(n19792) );
  nor2_1 U22696 ( .ip1(\pipeline/csr/mtime_full [10]), .ip2(n19792), .op(
        n19794) );
  nor3_1 U22697 ( .ip1(n21193), .ip2(n19794), .ip3(n20168), .op(n19793) );
  not_ab_or_c_or_d U22698 ( .ip1(n21195), .ip2(n19828), .ip3(n21120), .ip4(
        n19793), .op(n19797) );
  nor2_1 U22699 ( .ip1(n19794), .ip2(n20168), .op(n19795) );
  nor2_1 U22700 ( .ip1(n22254), .ip2(n19795), .op(n19796) );
  nor2_1 U22701 ( .ip1(n19797), .ip2(n19796), .op(\pipeline/csr/N2091 ) );
  nand2_1 U22702 ( .ip1(\pipeline/csr/mscratch [10]), .ip2(n22013), .op(n19799) );
  nand2_1 U22703 ( .ip1(n22014), .ip2(n19828), .op(n19798) );
  nand2_1 U22704 ( .ip1(n19799), .ip2(n19798), .op(n9918) );
  nand2_1 U22705 ( .ip1(\pipeline/csr/from_host [10]), .ip2(n22372), .op(
        n19801) );
  nand2_1 U22706 ( .ip1(n22373), .ip2(n19828), .op(n19800) );
  nand2_1 U22707 ( .ip1(n19801), .ip2(n19800), .op(n9950) );
  nand2_1 U22708 ( .ip1(n22378), .ip2(n19828), .op(n19803) );
  nand2_1 U22709 ( .ip1(\pipeline/csr/to_host [10]), .ip2(n22376), .op(n19802)
         );
  nand2_1 U22710 ( .ip1(n19803), .ip2(n19802), .op(n8762) );
  or2_1 U22711 ( .ip1(n19805), .ip2(n19804), .op(n19806) );
  nor2_1 U22712 ( .ip1(n21210), .ip2(n19806), .op(n19810) );
  not_ab_or_c_or_d U22713 ( .ip1(n19808), .ip2(n19807), .ip3(n22247), .ip4(
        n22157), .op(n19809) );
  or2_1 U22714 ( .ip1(n19810), .ip2(n19809), .op(\pipeline/csr/N2123 ) );
  or2_1 U22715 ( .ip1(\pipeline/csr/cycle_full [10]), .ip2(n19811), .op(n19812) );
  nand2_1 U22716 ( .ip1(n20187), .ip2(n19812), .op(n19813) );
  or2_1 U22717 ( .ip1(n21145), .ip2(n19813), .op(n19815) );
  nand2_1 U22718 ( .ip1(n22021), .ip2(n19828), .op(n19814) );
  nand2_1 U22719 ( .ip1(n19815), .ip2(n19814), .op(\pipeline/csr/N1883 ) );
  nand2_1 U22720 ( .ip1(\pipeline/csr/mtimecmp [10]), .ip2(n22363), .op(n19817) );
  nand2_1 U22721 ( .ip1(n22365), .ip2(n19828), .op(n19816) );
  nand2_1 U22722 ( .ip1(n19817), .ip2(n19816), .op(n10012) );
  mux2_1 U22723 ( .ip1(\pipeline/csr/instret_full [10]), .ip2(n19821), .s(
        n19818), .op(n19820) );
  nor2_1 U22724 ( .ip1(n21012), .ip2(n21011), .op(n19819) );
  nor2_1 U22725 ( .ip1(n19820), .ip2(n19819), .op(n19823) );
  nor2_1 U22726 ( .ip1(n19821), .ip2(n20990), .op(n19822) );
  nor2_1 U22727 ( .ip1(n19823), .ip2(n19822), .op(n19825) );
  nand2_1 U22728 ( .ip1(n21019), .ip2(n19828), .op(n19824) );
  nand2_1 U22729 ( .ip1(n19825), .ip2(n19824), .op(n10128) );
  nand2_1 U22730 ( .ip1(\pipeline/csr/mie [10]), .ip2(n22356), .op(n19827) );
  nand2_1 U22731 ( .ip1(n22357), .ip2(n19828), .op(n19826) );
  nand2_1 U22732 ( .ip1(n19827), .ip2(n19826), .op(n10050) );
  nand2_1 U22733 ( .ip1(n22314), .ip2(n19828), .op(n19832) );
  or2_1 U22734 ( .ip1(\pipeline/csr/cycle_full [42]), .ip2(n19829), .op(n19830) );
  nand3_1 U22735 ( .ip1(n20198), .ip2(n19830), .ip3(n22316), .op(n19831) );
  nand2_1 U22736 ( .ip1(n19832), .ip2(n19831), .op(\pipeline/csr/N1915 ) );
  inv_1 U22737 ( .ip(n19833), .op(n19834) );
  mux2_1 U22738 ( .ip1(\pipeline/csr_rdata_WB [10]), .ip2(n19834), .s(n17429), 
        .op(n8796) );
  nand2_1 U22739 ( .ip1(n21995), .ip2(imem_haddr[14]), .op(n19836) );
  nand2_1 U22740 ( .ip1(\pipeline/PC_IF [14]), .ip2(n21996), .op(n19835) );
  nand2_1 U22741 ( .ip1(n19836), .ip2(n19835), .op(n8462) );
  nand2_1 U22742 ( .ip1(\pipeline/PC_IF [14]), .ip2(n21988), .op(n19838) );
  nand2_1 U22743 ( .ip1(\pipeline/PC_DX [14]), .ip2(n21999), .op(n19837) );
  nand2_1 U22744 ( .ip1(n19838), .ip2(n19837), .op(n8461) );
  mux2_1 U22745 ( .ip1(\pipeline/PC_WB [14]), .ip2(\pipeline/PC_DX [14]), .s(
        n17777), .op(n8889) );
  nand2_1 U22746 ( .ip1(n21043), .ip2(n22171), .op(n19843) );
  xor2_1 U22747 ( .ip1(n19839), .ip2(\pipeline/PC_WB [14]), .op(n19840) );
  nand2_1 U22748 ( .ip1(n21046), .ip2(n19840), .op(n19842) );
  nand2_1 U22749 ( .ip1(\pipeline/epc [14]), .ip2(n21174), .op(n19841) );
  nand3_1 U22750 ( .ip1(n19843), .ip2(n19842), .ip3(n19841), .op(n8857) );
  nand2_1 U22751 ( .ip1(n21032), .ip2(n22171), .op(n19845) );
  nand2_1 U22752 ( .ip1(\pipeline/csr/mtvec [14]), .ip2(n20705), .op(n19844)
         );
  nand2_1 U22753 ( .ip1(n19845), .ip2(n19844), .op(n9978) );
  mux2_1 U22754 ( .ip1(dmem_haddr[14]), .ip2(\pipeline/alu_out_WB [14]), .s(
        n19505), .op(n8718) );
  nand2_1 U22755 ( .ip1(n22282), .ip2(n22171), .op(n19849) );
  or2_1 U22756 ( .ip1(\pipeline/csr/time_full [46]), .ip2(n20251), .op(n19846)
         );
  nand3_1 U22757 ( .ip1(n19847), .ip2(n19846), .ip3(n22284), .op(n19848) );
  nand2_1 U22758 ( .ip1(n19849), .ip2(n19848), .op(\pipeline/csr/N1983 ) );
  or2_1 U22759 ( .ip1(\pipeline/csr/time_full [14]), .ip2(n20246), .op(n19850)
         );
  nand2_1 U22760 ( .ip1(n19851), .ip2(n19850), .op(n19853) );
  nor2_1 U22761 ( .ip1(n21177), .ip2(n19853), .op(n19852) );
  not_ab_or_c_or_d U22762 ( .ip1(n21179), .ip2(n22171), .ip3(n21120), .ip4(
        n19852), .op(n19856) );
  inv_1 U22763 ( .ip(n19853), .op(n19854) );
  nor2_1 U22764 ( .ip1(n22254), .ip2(n19854), .op(n19855) );
  nor2_1 U22765 ( .ip1(n19856), .ip2(n19855), .op(\pipeline/csr/N1951 ) );
  inv_1 U22766 ( .ip(n19857), .op(n19858) );
  nor2_1 U22767 ( .ip1(\pipeline/csr/mtime_full [14]), .ip2(n19858), .op(
        n19861) );
  nor3_1 U22768 ( .ip1(n21193), .ip2(n19861), .ip3(n19860), .op(n19859) );
  not_ab_or_c_or_d U22769 ( .ip1(n21195), .ip2(n22171), .ip3(n21217), .ip4(
        n19859), .op(n19864) );
  nor2_1 U22770 ( .ip1(n19861), .ip2(n19860), .op(n19862) );
  nor2_1 U22771 ( .ip1(n22254), .ip2(n19862), .op(n19863) );
  nor2_1 U22772 ( .ip1(n19864), .ip2(n19863), .op(\pipeline/csr/N2095 ) );
  nand2_1 U22773 ( .ip1(\pipeline/csr/mscratch [14]), .ip2(n22013), .op(n19866) );
  nand2_1 U22774 ( .ip1(n22014), .ip2(n22171), .op(n19865) );
  nand2_1 U22775 ( .ip1(n19866), .ip2(n19865), .op(n9914) );
  nand2_1 U22776 ( .ip1(\pipeline/csr/from_host [14]), .ip2(n22372), .op(
        n19868) );
  nand2_1 U22777 ( .ip1(n22373), .ip2(n22171), .op(n19867) );
  nand2_1 U22778 ( .ip1(n19868), .ip2(n19867), .op(n9946) );
  nand2_1 U22779 ( .ip1(n22378), .ip2(n22171), .op(n19870) );
  nand2_1 U22780 ( .ip1(\pipeline/csr/to_host [14]), .ip2(n22376), .op(n19869)
         );
  nand2_1 U22781 ( .ip1(n19870), .ip2(n19869), .op(n8758) );
  or2_1 U22782 ( .ip1(\pipeline/csr/cycle_full [14]), .ip2(n20263), .op(n19871) );
  nand2_1 U22783 ( .ip1(n19872), .ip2(n19871), .op(n19873) );
  or2_1 U22784 ( .ip1(n21145), .ip2(n19873), .op(n19875) );
  nand2_1 U22785 ( .ip1(n22021), .ip2(n22171), .op(n19874) );
  nand2_1 U22786 ( .ip1(n19875), .ip2(n19874), .op(\pipeline/csr/N1887 ) );
  nand2_1 U22787 ( .ip1(\pipeline/csr/mtimecmp [14]), .ip2(n22363), .op(n19877) );
  nand2_1 U22788 ( .ip1(n22365), .ip2(n22171), .op(n19876) );
  nand2_1 U22789 ( .ip1(n19877), .ip2(n19876), .op(n10008) );
  mux2_1 U22790 ( .ip1(\pipeline/csr/instret_full [14]), .ip2(n19881), .s(
        n19878), .op(n19880) );
  nor2_1 U22791 ( .ip1(n21012), .ip2(n21011), .op(n19879) );
  nor2_1 U22792 ( .ip1(n19880), .ip2(n19879), .op(n19883) );
  nor2_1 U22793 ( .ip1(n19881), .ip2(n20990), .op(n19882) );
  nor2_1 U22794 ( .ip1(n19883), .ip2(n19882), .op(n19885) );
  nand2_1 U22795 ( .ip1(n21019), .ip2(n22171), .op(n19884) );
  nand2_1 U22796 ( .ip1(n19885), .ip2(n19884), .op(n10124) );
  nand2_1 U22797 ( .ip1(\pipeline/csr/mie [14]), .ip2(n22356), .op(n19887) );
  nand2_1 U22798 ( .ip1(n22357), .ip2(n22171), .op(n19886) );
  nand2_1 U22799 ( .ip1(n19887), .ip2(n19886), .op(n10046) );
  nand2_1 U22800 ( .ip1(n22314), .ip2(n22171), .op(n19891) );
  or2_1 U22801 ( .ip1(\pipeline/csr/cycle_full [46]), .ip2(n20271), .op(n19888) );
  nand3_1 U22802 ( .ip1(n19889), .ip2(n19888), .ip3(n22316), .op(n19890) );
  nand2_1 U22803 ( .ip1(n19891), .ip2(n19890), .op(\pipeline/csr/N1919 ) );
  mux2_1 U22804 ( .ip1(\pipeline/csr_rdata_WB [14]), .ip2(n19892), .s(n19498), 
        .op(n8792) );
  nor2_1 U22805 ( .ip1(n19894), .ip2(n10182), .op(n19895) );
  xor2_1 U22806 ( .ip1(n19896), .ip2(n19895), .op(imem_haddr[15]) );
  nand2_1 U22807 ( .ip1(n21995), .ip2(imem_haddr[15]), .op(n19898) );
  nand2_1 U22808 ( .ip1(\pipeline/PC_IF [15]), .ip2(n21996), .op(n19897) );
  nand2_1 U22809 ( .ip1(n19898), .ip2(n19897), .op(n8460) );
  nand2_1 U22810 ( .ip1(\pipeline/PC_IF [15]), .ip2(n21988), .op(n19900) );
  nand2_1 U22811 ( .ip1(\pipeline/PC_DX [15]), .ip2(n21999), .op(n19899) );
  nand2_1 U22812 ( .ip1(n19900), .ip2(n19899), .op(n8459) );
  mux2_1 U22813 ( .ip1(\pipeline/PC_WB [15]), .ip2(\pipeline/PC_DX [15]), .s(
        n17429), .op(n8888) );
  mux2_1 U22814 ( .ip1(\pipeline/PC_WB [16]), .ip2(\pipeline/PC_DX [16]), .s(
        n17777), .op(n8887) );
  inv_1 U22815 ( .ip(n19951), .op(n19901) );
  nor2_1 U22816 ( .ip1(n19901), .ip2(n21168), .op(n19906) );
  inv_1 U22817 ( .ip(\pipeline/PC_WB [16]), .op(n19904) );
  nand2_1 U22818 ( .ip1(n19902), .ip2(\pipeline/PC_WB [15]), .op(n19903) );
  not_ab_or_c_or_d U22819 ( .ip1(n19904), .ip2(n19903), .ip3(n19961), .ip4(
        n21171), .op(n19905) );
  ab_or_c_or_d U22820 ( .ip1(n21174), .ip2(\pipeline/epc [16]), .ip3(n19906), 
        .ip4(n19905), .op(n8855) );
  nand2_1 U22821 ( .ip1(n21032), .ip2(n19951), .op(n19908) );
  nand2_1 U22822 ( .ip1(\pipeline/csr/mtvec [16]), .ip2(n20705), .op(n19907)
         );
  nand2_1 U22823 ( .ip1(n19908), .ip2(n19907), .op(n9976) );
  mux2_1 U22824 ( .ip1(dmem_haddr[16]), .ip2(\pipeline/alu_out_WB [16]), .s(
        n21582), .op(n8716) );
  or2_1 U22825 ( .ip1(\pipeline/csr/time_full [16]), .ip2(n19909), .op(n19910)
         );
  nand2_1 U22826 ( .ip1(n19977), .ip2(n19910), .op(n19911) );
  or2_1 U22827 ( .ip1(n22002), .ip2(n19911), .op(n19913) );
  nand2_1 U22828 ( .ip1(n22005), .ip2(n19951), .op(n19912) );
  nand2_1 U22829 ( .ip1(n19913), .ip2(n19912), .op(\pipeline/csr/N1953 ) );
  inv_1 U22830 ( .ip(n19914), .op(n19915) );
  nor2_1 U22831 ( .ip1(\pipeline/csr/mtime_full [16]), .ip2(n19915), .op(
        n19917) );
  nor3_1 U22832 ( .ip1(n21193), .ip2(n19917), .ip3(n19966), .op(n19916) );
  not_ab_or_c_or_d U22833 ( .ip1(n21195), .ip2(n19951), .ip3(n21120), .ip4(
        n19916), .op(n19920) );
  nor2_1 U22834 ( .ip1(n19917), .ip2(n19966), .op(n19918) );
  nor2_1 U22835 ( .ip1(n21198), .ip2(n19918), .op(n19919) );
  nor2_1 U22836 ( .ip1(n19920), .ip2(n19919), .op(\pipeline/csr/N2097 ) );
  nand2_1 U22837 ( .ip1(\pipeline/csr/mscratch [16]), .ip2(n22013), .op(n19922) );
  nand2_1 U22838 ( .ip1(n22014), .ip2(n19951), .op(n19921) );
  nand2_1 U22839 ( .ip1(n19922), .ip2(n19921), .op(n9912) );
  nand2_1 U22840 ( .ip1(\pipeline/csr/from_host [16]), .ip2(n22372), .op(
        n19924) );
  nand2_1 U22841 ( .ip1(n22373), .ip2(n19951), .op(n19923) );
  nand2_1 U22842 ( .ip1(n19924), .ip2(n19923), .op(n9944) );
  nand2_1 U22843 ( .ip1(n22378), .ip2(n19951), .op(n19926) );
  nand2_1 U22844 ( .ip1(\pipeline/csr/to_host [16]), .ip2(n22376), .op(n19925)
         );
  nand2_1 U22845 ( .ip1(n19926), .ip2(n19925), .op(n8756) );
  or2_1 U22846 ( .ip1(n19927), .ip2(n22184), .op(n19929) );
  or2_1 U22847 ( .ip1(n22180), .ip2(n22184), .op(n19928) );
  nand2_1 U22848 ( .ip1(n19929), .ip2(n19928), .op(n19930) );
  nand2_1 U22849 ( .ip1(n18449), .ip2(n19930), .op(n19933) );
  nand2_1 U22850 ( .ip1(n21208), .ip2(n19951), .op(n19931) );
  or2_1 U22851 ( .ip1(n21210), .ip2(n19931), .op(n19932) );
  nand2_1 U22852 ( .ip1(n19933), .ip2(n19932), .op(\pipeline/csr/N2129 ) );
  or2_1 U22853 ( .ip1(\pipeline/csr/cycle_full [16]), .ip2(n19934), .op(n19935) );
  nand2_1 U22854 ( .ip1(n19985), .ip2(n19935), .op(n19936) );
  or2_1 U22855 ( .ip1(n21145), .ip2(n19936), .op(n19938) );
  nand2_1 U22856 ( .ip1(n22021), .ip2(n19951), .op(n19937) );
  nand2_1 U22857 ( .ip1(n19938), .ip2(n19937), .op(\pipeline/csr/N1889 ) );
  nand2_1 U22858 ( .ip1(\pipeline/csr/mtimecmp [16]), .ip2(n22363), .op(n19940) );
  nand2_1 U22859 ( .ip1(n22365), .ip2(n19951), .op(n19939) );
  nand2_1 U22860 ( .ip1(n19940), .ip2(n19939), .op(n10006) );
  mux2_1 U22861 ( .ip1(\pipeline/csr/instret_full [16]), .ip2(n19944), .s(
        n19941), .op(n19943) );
  nor2_1 U22862 ( .ip1(n21012), .ip2(n21011), .op(n19942) );
  nor2_1 U22863 ( .ip1(n19943), .ip2(n19942), .op(n19946) );
  nor2_1 U22864 ( .ip1(n19944), .ip2(n20990), .op(n19945) );
  nor2_1 U22865 ( .ip1(n19946), .ip2(n19945), .op(n19948) );
  nand2_1 U22866 ( .ip1(n21019), .ip2(n19951), .op(n19947) );
  nand2_1 U22867 ( .ip1(n19948), .ip2(n19947), .op(n10122) );
  nand2_1 U22868 ( .ip1(\pipeline/csr/mie [16]), .ip2(n22356), .op(n19950) );
  nand2_1 U22869 ( .ip1(n22357), .ip2(n19951), .op(n19949) );
  nand2_1 U22870 ( .ip1(n19950), .ip2(n19949), .op(n10044) );
  nand2_1 U22871 ( .ip1(n22314), .ip2(n19951), .op(n19955) );
  or2_1 U22872 ( .ip1(\pipeline/csr/cycle_full [48]), .ip2(n19952), .op(n19953) );
  nand3_1 U22873 ( .ip1(n20001), .ip2(n19953), .ip3(n22316), .op(n19954) );
  nand2_1 U22874 ( .ip1(n19955), .ip2(n19954), .op(\pipeline/csr/N1921 ) );
  mux2_1 U22875 ( .ip1(\pipeline/csr_rdata_WB [16]), .ip2(n19956), .s(n19498), 
        .op(n8790) );
  nand2_1 U22876 ( .ip1(n21995), .ip2(imem_haddr[17]), .op(n19958) );
  nand2_1 U22877 ( .ip1(\pipeline/PC_IF [17]), .ip2(n21996), .op(n19957) );
  nand2_1 U22878 ( .ip1(n19958), .ip2(n19957), .op(n8456) );
  nand2_1 U22879 ( .ip1(\pipeline/PC_IF [17]), .ip2(n22048), .op(n19960) );
  nand2_1 U22880 ( .ip1(\pipeline/PC_DX [17]), .ip2(n21999), .op(n19959) );
  nand2_1 U22881 ( .ip1(n19960), .ip2(n19959), .op(n8455) );
  mux2_1 U22882 ( .ip1(\pipeline/PC_WB [17]), .ip2(\pipeline/PC_DX [17]), .s(
        n17429), .op(n8886) );
  nand2_1 U22883 ( .ip1(n21043), .ip2(n22183), .op(n19965) );
  xor2_1 U22884 ( .ip1(n19961), .ip2(\pipeline/PC_WB [17]), .op(n19962) );
  nand2_1 U22885 ( .ip1(n21046), .ip2(n19962), .op(n19964) );
  nand2_1 U22886 ( .ip1(\pipeline/epc [17]), .ip2(n21174), .op(n19963) );
  nand3_1 U22887 ( .ip1(n19965), .ip2(n19964), .ip3(n19963), .op(n8854) );
  nand2_1 U22888 ( .ip1(n22008), .ip2(n22183), .op(n19969) );
  xor2_1 U22889 ( .ip1(n19966), .ip2(\pipeline/csr/mtime_full [17]), .op(
        n19967) );
  nand2_1 U22890 ( .ip1(n19967), .ip2(n22009), .op(n19968) );
  nand2_1 U22891 ( .ip1(n19969), .ip2(n19968), .op(\pipeline/csr/N2098 ) );
  nand2_1 U22892 ( .ip1(\pipeline/csr/mscratch [17]), .ip2(n22013), .op(n19971) );
  nand2_1 U22893 ( .ip1(n22014), .ip2(n22183), .op(n19970) );
  nand2_1 U22894 ( .ip1(n19971), .ip2(n19970), .op(n9911) );
  mux2_1 U22895 ( .ip1(dmem_haddr[17]), .ip2(\pipeline/alu_out_WB [17]), .s(
        n21582), .op(n8715) );
  inv_1 U22896 ( .ip(n22183), .op(n19998) );
  nor2_1 U22897 ( .ip1(n19998), .ip2(n22267), .op(n19976) );
  not_ab_or_c_or_d U22898 ( .ip1(n19974), .ip2(n19973), .ip3(n19972), .ip4(
        n22276), .op(n19975) );
  or2_1 U22899 ( .ip1(n19976), .ip2(n19975), .op(\pipeline/csr/N1986 ) );
  inv_1 U22900 ( .ip(n19977), .op(n19978) );
  nor2_1 U22901 ( .ip1(\pipeline/csr/time_full [17]), .ip2(n19978), .op(n19981) );
  nor3_1 U22902 ( .ip1(n21177), .ip2(n19980), .ip3(n19981), .op(n19979) );
  not_ab_or_c_or_d U22903 ( .ip1(n21179), .ip2(n22183), .ip3(n21217), .ip4(
        n19979), .op(n19984) );
  nor2_1 U22904 ( .ip1(n19981), .ip2(n19980), .op(n19982) );
  nor2_1 U22905 ( .ip1(n22254), .ip2(n19982), .op(n19983) );
  nor2_1 U22906 ( .ip1(n19984), .ip2(n19983), .op(\pipeline/csr/N1954 ) );
  inv_1 U22907 ( .ip(n19985), .op(n19986) );
  nor2_1 U22908 ( .ip1(\pipeline/csr/cycle_full [17]), .ip2(n19986), .op(
        n19989) );
  nor3_1 U22909 ( .ip1(n19988), .ip2(n19989), .ip3(n21215), .op(n19987) );
  not_ab_or_c_or_d U22910 ( .ip1(n21076), .ip2(n22183), .ip3(n21120), .ip4(
        n19987), .op(n19992) );
  nor2_1 U22911 ( .ip1(n19989), .ip2(n19988), .op(n19990) );
  nor2_1 U22912 ( .ip1(n21198), .ip2(n19990), .op(n19991) );
  nor2_1 U22913 ( .ip1(n19992), .ip2(n19991), .op(\pipeline/csr/N1890 ) );
  nor2_1 U22914 ( .ip1(n19998), .ip2(n21001), .op(n19997) );
  inv_1 U22915 ( .ip(\pipeline/csr/instret_full [17]), .op(n19994) );
  mux2_1 U22916 ( .ip1(n19994), .ip2(\pipeline/csr/instret_full [17]), .s(
        n19993), .op(n19995) );
  nor2_1 U22917 ( .ip1(n21005), .ip2(n19995), .op(n19996) );
  ab_or_c_or_d U22918 ( .ip1(n21016), .ip2(\pipeline/csr/instret_full [17]), 
        .ip3(n19997), .ip4(n19996), .op(n10121) );
  nor2_1 U22919 ( .ip1(n19998), .ip2(n22305), .op(n20003) );
  not_ab_or_c_or_d U22920 ( .ip1(n20001), .ip2(n20000), .ip3(n19999), .ip4(
        n22308), .op(n20002) );
  or2_1 U22921 ( .ip1(n20003), .ip2(n20002), .op(\pipeline/csr/N1922 ) );
  mux2_1 U22922 ( .ip1(\pipeline/csr_rdata_WB [17]), .ip2(n20004), .s(n17777), 
        .op(n8789) );
  nor2_1 U22923 ( .ip1(n20647), .ip2(n20005), .op(n20009) );
  nand2_1 U22924 ( .ip1(n20005), .ip2(n21649), .op(n20006) );
  nand2_1 U22925 ( .ip1(n20006), .ip2(n20649), .op(n20008) );
  mux2_1 U22926 ( .ip1(n20009), .ip2(n20008), .s(n20007), .op(n20016) );
  inv_1 U22927 ( .ip(n21643), .op(n21866) );
  xor2_1 U22928 ( .ip1(n20011), .ip2(n20010), .op(n20012) );
  nand2_1 U22929 ( .ip1(n14770), .ip2(n20012), .op(n20013) );
  xor2_1 U22930 ( .ip1(\pipeline/md/a [17]), .ip2(n20013), .op(n20014) );
  nor2_1 U22931 ( .ip1(n21866), .ip2(n20014), .op(n20015) );
  or2_1 U22932 ( .ip1(n20016), .ip2(n20015), .op(n8405) );
  inv_1 U22933 ( .ip(n20017), .op(n20018) );
  mux2_1 U22934 ( .ip1(\pipeline/csr_rdata_WB [18]), .ip2(n20018), .s(n19498), 
        .op(n8788) );
  inv_1 U22935 ( .ip(n20019), .op(n20020) );
  nor2_1 U22936 ( .ip1(n20021), .ip2(n20020), .op(n20022) );
  xor2_1 U22937 ( .ip1(n20022), .ip2(n20042), .op(imem_haddr[18]) );
  nand2_1 U22938 ( .ip1(n21995), .ip2(imem_haddr[18]), .op(n20024) );
  nand2_1 U22939 ( .ip1(\pipeline/PC_IF [18]), .ip2(n21996), .op(n20023) );
  nand2_1 U22940 ( .ip1(n20024), .ip2(n20023), .op(n8454) );
  nand2_1 U22941 ( .ip1(\pipeline/PC_IF [18]), .ip2(n21988), .op(n20026) );
  nand2_1 U22942 ( .ip1(\pipeline/PC_DX [18]), .ip2(n21999), .op(n20025) );
  nand2_1 U22943 ( .ip1(n20026), .ip2(n20025), .op(n8453) );
  mux2_1 U22944 ( .ip1(\pipeline/PC_WB [18]), .ip2(\pipeline/PC_DX [18]), .s(
        n17429), .op(n8885) );
  nor2_1 U22945 ( .ip1(n20027), .ip2(n21168), .op(n20034) );
  inv_1 U22946 ( .ip(\pipeline/PC_WB [19]), .op(n20032) );
  inv_1 U22947 ( .ip(n20028), .op(n20029) );
  nand2_1 U22948 ( .ip1(n20029), .ip2(\pipeline/PC_WB [18]), .op(n20031) );
  not_ab_or_c_or_d U22949 ( .ip1(n20032), .ip2(n20031), .ip3(n20030), .ip4(
        n21171), .op(n20033) );
  ab_or_c_or_d U22950 ( .ip1(n21174), .ip2(\pipeline/epc [19]), .ip3(n20034), 
        .ip4(n20033), .op(n8852) );
  nand2_1 U22951 ( .ip1(n20036), .ip2(n20035), .op(n20046) );
  xnor2_1 U22952 ( .ip1(n20046), .ip2(n20045), .op(imem_haddr[21]) );
  nand2_1 U22953 ( .ip1(n21995), .ip2(imem_haddr[21]), .op(n20048) );
  nand2_1 U22954 ( .ip1(\pipeline/PC_IF [21]), .ip2(n21996), .op(n20047) );
  nand2_1 U22955 ( .ip1(n20048), .ip2(n20047), .op(n8448) );
  nand2_1 U22956 ( .ip1(\pipeline/PC_IF [21]), .ip2(n22048), .op(n20050) );
  nand2_1 U22957 ( .ip1(\pipeline/PC_DX [21]), .ip2(n21999), .op(n20049) );
  nand2_1 U22958 ( .ip1(n20050), .ip2(n20049), .op(n8447) );
  mux2_1 U22959 ( .ip1(\pipeline/PC_WB [21]), .ip2(\pipeline/PC_DX [21]), .s(
        n17777), .op(n8882) );
  mux2_1 U22960 ( .ip1(\pipeline/PC_WB [22]), .ip2(\pipeline/PC_DX [22]), .s(
        n19498), .op(n8881) );
  nor2_1 U22961 ( .ip1(n22203), .ip2(n21168), .op(n20056) );
  inv_1 U22962 ( .ip(\pipeline/PC_WB [22]), .op(n20054) );
  inv_1 U22963 ( .ip(n20051), .op(n20052) );
  nand2_1 U22964 ( .ip1(n20052), .ip2(\pipeline/PC_WB [21]), .op(n20053) );
  not_ab_or_c_or_d U22965 ( .ip1(n20054), .ip2(n20053), .ip3(n20110), .ip4(
        n21171), .op(n20055) );
  ab_or_c_or_d U22966 ( .ip1(n21174), .ip2(\pipeline/epc [22]), .ip3(n20056), 
        .ip4(n20055), .op(n8849) );
  nand2_1 U22967 ( .ip1(n21032), .ip2(n20100), .op(n20058) );
  nand2_1 U22968 ( .ip1(\pipeline/csr/mtvec [22]), .ip2(n20705), .op(n20057)
         );
  nand2_1 U22969 ( .ip1(n20058), .ip2(n20057), .op(n9970) );
  mux2_1 U22970 ( .ip1(dmem_haddr[22]), .ip2(\pipeline/alu_out_WB [22]), .s(
        n21582), .op(n8710) );
  nand2_1 U22971 ( .ip1(n22282), .ip2(n20100), .op(n20062) );
  or2_1 U22972 ( .ip1(\pipeline/csr/time_full [54]), .ip2(n20059), .op(n20060)
         );
  nand3_1 U22973 ( .ip1(n20060), .ip2(n22277), .ip3(n22284), .op(n20061) );
  nand2_1 U22974 ( .ip1(n20062), .ip2(n20061), .op(\pipeline/csr/N1991 ) );
  or2_1 U22975 ( .ip1(\pipeline/csr/time_full [22]), .ip2(n20063), .op(n20064)
         );
  nand2_1 U22976 ( .ip1(n20115), .ip2(n20064), .op(n20066) );
  nor2_1 U22977 ( .ip1(n21177), .ip2(n20066), .op(n20065) );
  not_ab_or_c_or_d U22978 ( .ip1(n21179), .ip2(n20100), .ip3(n21217), .ip4(
        n20065), .op(n20069) );
  inv_1 U22979 ( .ip(n20066), .op(n20067) );
  nor2_1 U22980 ( .ip1(n21198), .ip2(n20067), .op(n20068) );
  nor2_1 U22981 ( .ip1(n20069), .ip2(n20068), .op(\pipeline/csr/N1959 ) );
  inv_1 U22982 ( .ip(n20070), .op(n20071) );
  nor2_1 U22983 ( .ip1(\pipeline/csr/mtime_full [22]), .ip2(n20071), .op(
        n20073) );
  nor3_1 U22984 ( .ip1(n21193), .ip2(n20073), .ip3(n20123), .op(n20072) );
  not_ab_or_c_or_d U22985 ( .ip1(n21195), .ip2(n20100), .ip3(n21120), .ip4(
        n20072), .op(n20076) );
  nor2_1 U22986 ( .ip1(n20073), .ip2(n20123), .op(n20074) );
  nor2_1 U22987 ( .ip1(n22254), .ip2(n20074), .op(n20075) );
  nor2_1 U22988 ( .ip1(n20076), .ip2(n20075), .op(\pipeline/csr/N2103 ) );
  nand2_1 U22989 ( .ip1(\pipeline/csr/mscratch [22]), .ip2(n22013), .op(n20078) );
  nand2_1 U22990 ( .ip1(n22014), .ip2(n20100), .op(n20077) );
  nand2_1 U22991 ( .ip1(n20078), .ip2(n20077), .op(n9906) );
  nand2_1 U22992 ( .ip1(\pipeline/csr/from_host [22]), .ip2(n22372), .op(
        n20080) );
  nand2_1 U22993 ( .ip1(n22373), .ip2(n20100), .op(n20079) );
  nand2_1 U22994 ( .ip1(n20080), .ip2(n20079), .op(n9938) );
  nand2_1 U22995 ( .ip1(n22378), .ip2(n20100), .op(n20082) );
  nand2_1 U22996 ( .ip1(\pipeline/csr/to_host [22]), .ip2(n22376), .op(n20081)
         );
  nand2_1 U22997 ( .ip1(n20082), .ip2(n20081), .op(n8750) );
  or2_1 U22998 ( .ip1(\pipeline/csr/cycle_full [22]), .ip2(n20083), .op(n20084) );
  nand2_1 U22999 ( .ip1(n20133), .ip2(n20084), .op(n20085) );
  or2_1 U23000 ( .ip1(n21145), .ip2(n20085), .op(n20087) );
  nand2_1 U23001 ( .ip1(n22021), .ip2(n20100), .op(n20086) );
  nand2_1 U23002 ( .ip1(n20087), .ip2(n20086), .op(\pipeline/csr/N1895 ) );
  nand2_1 U23003 ( .ip1(\pipeline/csr/mtimecmp [22]), .ip2(n22363), .op(n20089) );
  nand2_1 U23004 ( .ip1(n22365), .ip2(n20100), .op(n20088) );
  nand2_1 U23005 ( .ip1(n20089), .ip2(n20088), .op(n10000) );
  mux2_1 U23006 ( .ip1(\pipeline/csr/instret_full [22]), .ip2(n20093), .s(
        n20090), .op(n20092) );
  nor2_1 U23007 ( .ip1(n21012), .ip2(n21011), .op(n20091) );
  nor2_1 U23008 ( .ip1(n20092), .ip2(n20091), .op(n20095) );
  nor2_1 U23009 ( .ip1(n20093), .ip2(n20990), .op(n20094) );
  nor2_1 U23010 ( .ip1(n20095), .ip2(n20094), .op(n20097) );
  nand2_1 U23011 ( .ip1(n21019), .ip2(n20100), .op(n20096) );
  nand2_1 U23012 ( .ip1(n20097), .ip2(n20096), .op(n10116) );
  nand2_1 U23013 ( .ip1(\pipeline/csr/mie [22]), .ip2(n22356), .op(n20099) );
  nand2_1 U23014 ( .ip1(n22357), .ip2(n20100), .op(n20098) );
  nand2_1 U23015 ( .ip1(n20099), .ip2(n20098), .op(n10038) );
  nand2_1 U23016 ( .ip1(n22314), .ip2(n20100), .op(n20104) );
  or2_1 U23017 ( .ip1(\pipeline/csr/cycle_full [54]), .ip2(n20101), .op(n20102) );
  nand3_1 U23018 ( .ip1(n20102), .ip2(n22301), .ip3(n22316), .op(n20103) );
  nand2_1 U23019 ( .ip1(n20104), .ip2(n20103), .op(\pipeline/csr/N1927 ) );
  mux2_1 U23020 ( .ip1(\pipeline/csr_rdata_WB [22]), .ip2(n20105), .s(n20389), 
        .op(n8784) );
  nand2_1 U23021 ( .ip1(\pipeline/PC_IF [23]), .ip2(n21996), .op(n20106) );
  nand2_1 U23022 ( .ip1(n20107), .ip2(n20106), .op(n8444) );
  nand2_1 U23023 ( .ip1(\pipeline/PC_IF [23]), .ip2(n21988), .op(n20109) );
  nand2_1 U23024 ( .ip1(\pipeline/PC_DX [23]), .ip2(n21999), .op(n20108) );
  nand2_1 U23025 ( .ip1(n20109), .ip2(n20108), .op(n8443) );
  mux2_1 U23026 ( .ip1(\pipeline/PC_WB [23]), .ip2(\pipeline/PC_DX [23]), .s(
        n20389), .op(n8880) );
  nand2_1 U23027 ( .ip1(n21043), .ip2(n22274), .op(n20114) );
  xor2_1 U23028 ( .ip1(n20110), .ip2(\pipeline/PC_WB [23]), .op(n20111) );
  nand2_1 U23029 ( .ip1(n21046), .ip2(n20111), .op(n20113) );
  nand2_1 U23030 ( .ip1(\pipeline/epc [23]), .ip2(n21174), .op(n20112) );
  nand3_1 U23031 ( .ip1(n20114), .ip2(n20113), .ip3(n20112), .op(n8848) );
  mux2_1 U23032 ( .ip1(dmem_haddr[23]), .ip2(\pipeline/alu_out_WB [23]), .s(
        n21582), .op(n8709) );
  inv_1 U23033 ( .ip(n20115), .op(n20116) );
  nor2_1 U23034 ( .ip1(\pipeline/csr/time_full [23]), .ip2(n20116), .op(n20119) );
  nor3_1 U23035 ( .ip1(n21177), .ip2(n20118), .ip3(n20119), .op(n20117) );
  not_ab_or_c_or_d U23036 ( .ip1(n21179), .ip2(n22274), .ip3(n21217), .ip4(
        n20117), .op(n20122) );
  nor2_1 U23037 ( .ip1(n20119), .ip2(n20118), .op(n20120) );
  nor2_1 U23038 ( .ip1(n22254), .ip2(n20120), .op(n20121) );
  nor2_1 U23039 ( .ip1(n20122), .ip2(n20121), .op(\pipeline/csr/N1960 ) );
  nand2_1 U23040 ( .ip1(n22008), .ip2(n22274), .op(n20126) );
  xor2_1 U23041 ( .ip1(n20123), .ip2(\pipeline/csr/mtime_full [23]), .op(
        n20124) );
  nand2_1 U23042 ( .ip1(n20124), .ip2(n22009), .op(n20125) );
  nand2_1 U23043 ( .ip1(n20126), .ip2(n20125), .op(\pipeline/csr/N2104 ) );
  nand2_1 U23044 ( .ip1(\pipeline/csr/mscratch [23]), .ip2(n22013), .op(n20128) );
  nand2_1 U23045 ( .ip1(n22014), .ip2(n22274), .op(n20127) );
  nand2_1 U23046 ( .ip1(n20128), .ip2(n20127), .op(n9905) );
  nand2_1 U23047 ( .ip1(\pipeline/csr/from_host [23]), .ip2(n22372), .op(
        n20130) );
  nand2_1 U23048 ( .ip1(n22373), .ip2(n22274), .op(n20129) );
  nand2_1 U23049 ( .ip1(n20130), .ip2(n20129), .op(n9937) );
  nand2_1 U23050 ( .ip1(n22378), .ip2(n22274), .op(n20132) );
  nand2_1 U23051 ( .ip1(\pipeline/csr/to_host [23]), .ip2(n22376), .op(n20131)
         );
  nand2_1 U23052 ( .ip1(n20132), .ip2(n20131), .op(n8749) );
  inv_1 U23053 ( .ip(n20133), .op(n20134) );
  nor2_1 U23054 ( .ip1(\pipeline/csr/cycle_full [23]), .ip2(n20134), .op(
        n20137) );
  nor3_1 U23055 ( .ip1(n20136), .ip2(n20137), .ip3(n21215), .op(n20135) );
  not_ab_or_c_or_d U23056 ( .ip1(n21076), .ip2(n22274), .ip3(n21120), .ip4(
        n20135), .op(n20140) );
  nor2_1 U23057 ( .ip1(n20137), .ip2(n20136), .op(n20138) );
  nor2_1 U23058 ( .ip1(n21198), .ip2(n20138), .op(n20139) );
  nor2_1 U23059 ( .ip1(n20140), .ip2(n20139), .op(\pipeline/csr/N1896 ) );
  nand2_1 U23060 ( .ip1(\pipeline/csr/mtimecmp [23]), .ip2(n22363), .op(n20142) );
  nand2_1 U23061 ( .ip1(n22365), .ip2(n22274), .op(n20141) );
  nand2_1 U23062 ( .ip1(n20142), .ip2(n20141), .op(n9999) );
  nand2_1 U23063 ( .ip1(\pipeline/csr/mie [23]), .ip2(n22356), .op(n20144) );
  nand2_1 U23064 ( .ip1(n22357), .ip2(n22274), .op(n20143) );
  nand2_1 U23065 ( .ip1(n20144), .ip2(n20143), .op(n10037) );
  mux2_1 U23066 ( .ip1(\pipeline/csr_rdata_WB [23]), .ip2(n20145), .s(n20389), 
        .op(n8783) );
  inv_1 U23067 ( .ip(n20149), .op(n20147) );
  inv_1 U23068 ( .ip(n21944), .op(n21730) );
  nor3_1 U23069 ( .ip1(n20147), .ip2(n20146), .ip3(n21730), .op(n20156) );
  nor2_1 U23070 ( .ip1(n20149), .ip2(n20148), .op(n20153) );
  nor2_1 U23071 ( .ip1(n20151), .ip2(n20150), .op(n20152) );
  nor2_1 U23072 ( .ip1(n20153), .ip2(n20152), .op(n20154) );
  nor2_1 U23073 ( .ip1(n20154), .ip2(n22665), .op(n20155) );
  not_ab_or_c_or_d U23074 ( .ip1(n21884), .ip2(\pipeline/md/a [25]), .ip3(
        n20156), .ip4(n20155), .op(n20161) );
  xor2_1 U23075 ( .ip1(n20158), .ip2(n20157), .op(n20159) );
  nand2_1 U23076 ( .ip1(n21649), .ip2(n20159), .op(n20160) );
  nand2_1 U23077 ( .ip1(n20161), .ip2(n20160), .op(n8397) );
  mux2_1 U23078 ( .ip1(\pipeline/csr_rdata_WB [25]), .ip2(n20162), .s(n20389), 
        .op(n8781) );
  mux2_1 U23079 ( .ip1(\pipeline/csr_rdata_WB [27]), .ip2(n20163), .s(n20389), 
        .op(n8779) );
  nand2_1 U23080 ( .ip1(n21995), .ip2(imem_haddr[28]), .op(n20165) );
  nand2_1 U23081 ( .ip1(\pipeline/PC_IF [28]), .ip2(n21996), .op(n20164) );
  nand2_1 U23082 ( .ip1(n20165), .ip2(n20164), .op(n8434) );
  nand2_1 U23083 ( .ip1(\pipeline/PC_IF [28]), .ip2(n21988), .op(n20167) );
  nand2_1 U23084 ( .ip1(\pipeline/PC_DX [28]), .ip2(n21999), .op(n20166) );
  nand2_1 U23085 ( .ip1(n20167), .ip2(n20166), .op(n8433) );
  mux2_1 U23086 ( .ip1(dmem_haddr[11]), .ip2(\pipeline/alu_out_WB [11]), .s(
        n19505), .op(n8721) );
  nand2_1 U23087 ( .ip1(n22008), .ip2(n22156), .op(n20171) );
  xor2_1 U23088 ( .ip1(n20168), .ip2(\pipeline/csr/mtime_full [11]), .op(
        n20169) );
  nand2_1 U23089 ( .ip1(n20169), .ip2(n22009), .op(n20170) );
  nand2_1 U23090 ( .ip1(n20171), .ip2(n20170), .op(\pipeline/csr/N2092 ) );
  nand2_1 U23091 ( .ip1(\pipeline/csr/mscratch [11]), .ip2(n22013), .op(n20173) );
  nand2_1 U23092 ( .ip1(n22014), .ip2(n22156), .op(n20172) );
  nand2_1 U23093 ( .ip1(n20173), .ip2(n20172), .op(n9917) );
  nor2_1 U23094 ( .ip1(n20196), .ip2(n22267), .op(n20177) );
  not_ab_or_c_or_d U23095 ( .ip1(n20175), .ip2(n20174), .ip3(n22276), .ip4(
        n20747), .op(n20176) );
  or2_1 U23096 ( .ip1(n20177), .ip2(n20176), .op(\pipeline/csr/N1980 ) );
  inv_1 U23097 ( .ip(n20183), .op(n20178) );
  nor2_1 U23098 ( .ip1(\pipeline/csr/time_full [11]), .ip2(n20178), .op(n20179) );
  nor2_1 U23099 ( .ip1(n20752), .ip2(n20179), .op(n20180) );
  nor2_1 U23100 ( .ip1(n22254), .ip2(n20180), .op(n20182) );
  inv_1 U23101 ( .ip(n20181), .op(n22255) );
  not_ab_or_c_or_d U23102 ( .ip1(n20196), .ip2(n22257), .ip3(n20182), .ip4(
        n22255), .op(n20186) );
  not_ab_or_c_or_d U23103 ( .ip1(n20184), .ip2(n20183), .ip3(n21177), .ip4(
        n20752), .op(n20185) );
  or2_1 U23104 ( .ip1(n20186), .ip2(n20185), .op(\pipeline/csr/N1948 ) );
  inv_1 U23105 ( .ip(n20187), .op(n20188) );
  nor2_1 U23106 ( .ip1(\pipeline/csr/cycle_full [11]), .ip2(n20188), .op(
        n20190) );
  nor3_1 U23107 ( .ip1(n20772), .ip2(n20190), .ip3(n21215), .op(n20189) );
  not_ab_or_c_or_d U23108 ( .ip1(n21076), .ip2(n22156), .ip3(n21217), .ip4(
        n20189), .op(n20193) );
  nor2_1 U23109 ( .ip1(n20190), .ip2(n20772), .op(n20191) );
  nor2_1 U23110 ( .ip1(n22254), .ip2(n20191), .op(n20192) );
  nor2_1 U23111 ( .ip1(n20193), .ip2(n20192), .op(\pipeline/csr/N1884 ) );
  nand2_1 U23112 ( .ip1(\pipeline/csr/mie [11]), .ip2(n22356), .op(n20195) );
  nand2_1 U23113 ( .ip1(n22357), .ip2(n22156), .op(n20194) );
  nand2_1 U23114 ( .ip1(n20195), .ip2(n20194), .op(n10049) );
  nor2_1 U23115 ( .ip1(n20196), .ip2(n22305), .op(n20200) );
  not_ab_or_c_or_d U23116 ( .ip1(n20198), .ip2(n20197), .ip3(n22308), .ip4(
        n20789), .op(n20199) );
  or2_1 U23117 ( .ip1(n20200), .ip2(n20199), .op(\pipeline/csr/N1916 ) );
  inv_1 U23118 ( .ip(n20201), .op(n20202) );
  mux2_1 U23119 ( .ip1(\pipeline/csr_rdata_WB [11]), .ip2(n20202), .s(n20389), 
        .op(n8795) );
  nand2_1 U23120 ( .ip1(imem_haddr[13]), .ip2(n21995), .op(n20204) );
  nand2_1 U23121 ( .ip1(\pipeline/PC_IF [13]), .ip2(n21996), .op(n20203) );
  nand2_1 U23122 ( .ip1(n20204), .ip2(n20203), .op(n8464) );
  nand2_1 U23123 ( .ip1(\pipeline/PC_IF [13]), .ip2(n21988), .op(n20206) );
  nand2_1 U23124 ( .ip1(\pipeline/PC_DX [13]), .ip2(n21999), .op(n20205) );
  nand2_1 U23125 ( .ip1(n20206), .ip2(n20205), .op(n8463) );
  mux2_1 U23126 ( .ip1(\pipeline/PC_WB [13]), .ip2(\pipeline/PC_DX [13]), .s(
        n20389), .op(n8890) );
  nand2_1 U23127 ( .ip1(n20208), .ip2(n20207), .op(n20214) );
  nand2_1 U23128 ( .ip1(n20210), .ip2(n20209), .op(n20211) );
  nand2_1 U23129 ( .ip1(n20212), .ip2(n20211), .op(n20213) );
  xnor2_1 U23130 ( .ip1(n20214), .ip2(n20213), .op(n20215) );
  nand2_1 U23131 ( .ip1(n20215), .ip2(n21577), .op(n20243) );
  inv_1 U23132 ( .ip(n20216), .op(n20217) );
  nor2_1 U23133 ( .ip1(n20726), .ip2(n20217), .op(n20237) );
  or2_1 U23134 ( .ip1(n20219), .ip2(n20218), .op(n20235) );
  nor3_1 U23135 ( .ip1(n20220), .ip2(n21551), .ip3(n13678), .op(n20225) );
  nor2_1 U23136 ( .ip1(n20222), .ip2(n20221), .op(n20223) );
  nor2_1 U23137 ( .ip1(n20907), .ip2(n20223), .op(n20224) );
  not_ab_or_c_or_d U23138 ( .ip1(n20911), .ip2(n20226), .ip3(n20225), .ip4(
        n20224), .op(n20234) );
  inv_1 U23139 ( .ip(n20227), .op(n20228) );
  nand2_1 U23140 ( .ip1(n20229), .ip2(n20228), .op(n20233) );
  nand2_1 U23141 ( .ip1(n20231), .ip2(n20230), .op(n20232) );
  not_ab_or_c_or_d U23142 ( .ip1(n20239), .ip2(n20238), .ip3(n20237), .ip4(
        n20236), .op(n20242) );
  nand2_1 U23143 ( .ip1(n20240), .ip2(n20900), .op(n20241) );
  nand3_1 U23144 ( .ip1(n20243), .ip2(n20242), .ip3(n20241), .op(
        dmem_haddr[13]) );
  mux2_1 U23145 ( .ip1(dmem_haddr[13]), .ip2(\pipeline/alu_out_WB [13]), .s(
        n21582), .op(n8719) );
  inv_1 U23146 ( .ip(n20754), .op(n20244) );
  nor2_1 U23147 ( .ip1(\pipeline/csr/time_full [13]), .ip2(n20244), .op(n20247) );
  nor3_1 U23148 ( .ip1(n21177), .ip2(n20246), .ip3(n20247), .op(n20245) );
  not_ab_or_c_or_d U23149 ( .ip1(n21179), .ip2(n22166), .ip3(n21120), .ip4(
        n20245), .op(n20250) );
  nor2_1 U23150 ( .ip1(n20247), .ip2(n20246), .op(n20248) );
  nor2_1 U23151 ( .ip1(n21198), .ip2(n20248), .op(n20249) );
  nor2_1 U23152 ( .ip1(n20250), .ip2(n20249), .op(\pipeline/csr/N1950 ) );
  nor2_1 U23153 ( .ip1(n20270), .ip2(n22267), .op(n20255) );
  not_ab_or_c_or_d U23154 ( .ip1(n20253), .ip2(n20252), .ip3(n20251), .ip4(
        n22276), .op(n20254) );
  or2_1 U23155 ( .ip1(n20255), .ip2(n20254), .op(\pipeline/csr/N1982 ) );
  nand2_1 U23156 ( .ip1(n22008), .ip2(n22166), .op(n20258) );
  xor2_1 U23157 ( .ip1(\pipeline/csr/mtime_full [13]), .ip2(n20761), .op(
        n20256) );
  nand2_1 U23158 ( .ip1(n20256), .ip2(n22009), .op(n20257) );
  nand2_1 U23159 ( .ip1(n20258), .ip2(n20257), .op(\pipeline/csr/N2094 ) );
  nand2_1 U23160 ( .ip1(\pipeline/csr/mscratch [13]), .ip2(n22013), .op(n20260) );
  nand2_1 U23161 ( .ip1(n22014), .ip2(n22166), .op(n20259) );
  nand2_1 U23162 ( .ip1(n20260), .ip2(n20259), .op(n9915) );
  inv_1 U23163 ( .ip(n20774), .op(n20261) );
  nor2_1 U23164 ( .ip1(\pipeline/csr/cycle_full [13]), .ip2(n20261), .op(
        n20264) );
  nor3_1 U23165 ( .ip1(n20263), .ip2(n20264), .ip3(n21215), .op(n20262) );
  not_ab_or_c_or_d U23166 ( .ip1(n21076), .ip2(n22166), .ip3(n21217), .ip4(
        n20262), .op(n20267) );
  nor2_1 U23167 ( .ip1(n20264), .ip2(n20263), .op(n20265) );
  nor2_1 U23168 ( .ip1(n21198), .ip2(n20265), .op(n20266) );
  nor2_1 U23169 ( .ip1(n20267), .ip2(n20266), .op(\pipeline/csr/N1886 ) );
  nand2_1 U23170 ( .ip1(\pipeline/csr/mie [13]), .ip2(n22356), .op(n20269) );
  nand2_1 U23171 ( .ip1(n22357), .ip2(n22166), .op(n20268) );
  nand2_1 U23172 ( .ip1(n20269), .ip2(n20268), .op(n10047) );
  nor2_1 U23173 ( .ip1(n20270), .ip2(n22305), .op(n20274) );
  not_ab_or_c_or_d U23174 ( .ip1(n20791), .ip2(n20272), .ip3(n20271), .ip4(
        n22308), .op(n20273) );
  or2_1 U23175 ( .ip1(n20274), .ip2(n20273), .op(\pipeline/csr/N1918 ) );
  mux2_1 U23176 ( .ip1(\pipeline/csr_rdata_WB [13]), .ip2(n20275), .s(n20389), 
        .op(n8793) );
  nand2_1 U23177 ( .ip1(n21649), .ip2(n20277), .op(n20276) );
  nand2_1 U23178 ( .ip1(n20649), .ip2(n20276), .op(n20280) );
  nor2_1 U23179 ( .ip1(n20277), .ip2(n20647), .op(n20279) );
  mux2_1 U23180 ( .ip1(n20280), .ip2(n20279), .s(n20278), .op(n20291) );
  nor2_1 U23181 ( .ip1(n20282), .ip2(n20281), .op(n20603) );
  nor2_1 U23182 ( .ip1(n20283), .ip2(n20603), .op(n20284) );
  nor2_1 U23183 ( .ip1(n20285), .ip2(n20284), .op(n20286) );
  xor2_1 U23184 ( .ip1(\pipeline/md/b [23]), .ip2(n20286), .op(n20287) );
  nand2_1 U23185 ( .ip1(n20287), .ip2(n14770), .op(n20288) );
  xor2_1 U23186 ( .ip1(\pipeline/md/a [23]), .ip2(n20288), .op(n20289) );
  nor2_1 U23187 ( .ip1(n21866), .ip2(n20289), .op(n20290) );
  or2_1 U23188 ( .ip1(n20291), .ip2(n20290), .op(n8408) );
  nor4_1 U23189 ( .ip1(\pipeline/md_resp_result [26]), .ip2(n20308), .ip3(
        n20307), .ip4(n22755), .op(n20305) );
  nand2_1 U23190 ( .ip1(\pipeline/md/negate_output ), .ip2(n20292), .op(n20294) );
  nor2_1 U23191 ( .ip1(n20295), .ip2(n20294), .op(n20293) );
  not_ab_or_c_or_d U23192 ( .ip1(n20295), .ip2(n20294), .ip3(n21960), .ip4(
        n20293), .op(n20303) );
  nand2_1 U23193 ( .ip1(\pipeline/md/negate_output ), .ip2(n20296), .op(n20297) );
  nor2_1 U23194 ( .ip1(\pipeline/md/result [58]), .ip2(n20297), .op(n20299) );
  and2_1 U23195 ( .ip1(\pipeline/md/result [58]), .ip2(n20297), .op(n20298) );
  nor2_1 U23196 ( .ip1(n20299), .ip2(n20298), .op(n20300) );
  nor2_1 U23197 ( .ip1(n20300), .ip2(n21967), .op(n20301) );
  nor2_1 U23198 ( .ip1(n21972), .ip2(n20301), .op(n20302) );
  nor2_1 U23199 ( .ip1(n20303), .ip2(n20302), .op(n20304) );
  not_ab_or_c_or_d U23200 ( .ip1(n21978), .ip2(n20306), .ip3(n20305), .ip4(
        n20304), .op(n20314) );
  or2_1 U23201 ( .ip1(n20308), .ip2(n20307), .op(n20309) );
  nand2_1 U23202 ( .ip1(n20310), .ip2(n20309), .op(n20311) );
  nand2_1 U23203 ( .ip1(n22738), .ip2(n20311), .op(n20312) );
  nand2_1 U23204 ( .ip1(\pipeline/md_resp_result [26]), .ip2(n20312), .op(
        n20313) );
  nand2_1 U23205 ( .ip1(n20314), .ip2(n20313), .op(n8608) );
  mux2_1 U23206 ( .ip1(\pipeline/csr_rdata_WB [26]), .ip2(n20315), .s(n20389), 
        .op(n8780) );
  nand2_1 U23207 ( .ip1(imem_haddr[29]), .ip2(n21995), .op(n20317) );
  nand2_1 U23208 ( .ip1(\pipeline/PC_IF [29]), .ip2(n21996), .op(n20316) );
  nand2_1 U23209 ( .ip1(n20317), .ip2(n20316), .op(n8432) );
  nand2_1 U23210 ( .ip1(\pipeline/PC_IF [29]), .ip2(n21988), .op(n20319) );
  nand2_1 U23211 ( .ip1(\pipeline/PC_DX [29]), .ip2(n21999), .op(n20318) );
  nand2_1 U23212 ( .ip1(n20319), .ip2(n20318), .op(n8431) );
  mux2_1 U23213 ( .ip1(\pipeline/PC_WB [29]), .ip2(\pipeline/PC_DX [29]), .s(
        n20389), .op(n8874) );
  nand2_1 U23214 ( .ip1(n21043), .ip2(n22234), .op(n20324) );
  xor2_1 U23215 ( .ip1(n20320), .ip2(\pipeline/PC_WB [29]), .op(n20321) );
  nand2_1 U23216 ( .ip1(n21046), .ip2(n20321), .op(n20323) );
  nand2_1 U23217 ( .ip1(\pipeline/epc [29]), .ip2(n21174), .op(n20322) );
  nand3_1 U23218 ( .ip1(n20324), .ip2(n20323), .ip3(n20322), .op(n8842) );
  nand2_1 U23219 ( .ip1(n21995), .ip2(imem_haddr[30]), .op(n20326) );
  nand2_1 U23220 ( .ip1(\pipeline/PC_IF [30]), .ip2(n21996), .op(n20325) );
  nand2_1 U23221 ( .ip1(n20326), .ip2(n20325), .op(n8430) );
  nand2_1 U23222 ( .ip1(\pipeline/PC_IF [30]), .ip2(n21988), .op(n20328) );
  nand2_1 U23223 ( .ip1(\pipeline/PC_DX [30]), .ip2(n21999), .op(n20327) );
  nand2_1 U23224 ( .ip1(n20328), .ip2(n20327), .op(n8429) );
  mux2_1 U23225 ( .ip1(dmem_haddr[6]), .ip2(\pipeline/alu_out_WB [6]), .s(
        n19505), .op(n8726) );
  nand2_1 U23226 ( .ip1(n22282), .ip2(n22364), .op(n20332) );
  or2_1 U23227 ( .ip1(\pipeline/csr/time_full [38]), .ip2(n21050), .op(n20329)
         );
  nand3_1 U23228 ( .ip1(n20330), .ip2(n20329), .ip3(n22284), .op(n20331) );
  nand2_1 U23229 ( .ip1(n20332), .ip2(n20331), .op(\pipeline/csr/N1975 ) );
  nand2_1 U23230 ( .ip1(n20844), .ip2(n22145), .op(n20337) );
  nand2_1 U23231 ( .ip1(n21117), .ip2(\pipeline/csr/instret_full [37]), .op(
        n20336) );
  or2_1 U23232 ( .ip1(\pipeline/csr/instret_full [37]), .ip2(n20809), .op(
        n20333) );
  nand3_1 U23233 ( .ip1(n20334), .ip2(n20340), .ip3(n20333), .op(n20335) );
  nand3_1 U23234 ( .ip1(n20337), .ip2(n20336), .ip3(n20335), .op(n10101) );
  nor2_1 U23235 ( .ip1(n19134), .ip2(n20339), .op(n20342) );
  not_ab_or_c_or_d U23236 ( .ip1(n20340), .ip2(n20339), .ip3(n20338), .ip4(
        n21111), .op(n20341) );
  ab_or_c_or_d U23237 ( .ip1(n20844), .ip2(n22364), .ip3(n20342), .ip4(n20341), 
        .op(n10100) );
  or2_1 U23238 ( .ip1(\pipeline/csr/time_full [6]), .ip2(n21058), .op(n20343)
         );
  nand2_1 U23239 ( .ip1(n20344), .ip2(n20343), .op(n20346) );
  nor2_1 U23240 ( .ip1(n21177), .ip2(n20346), .op(n20345) );
  not_ab_or_c_or_d U23241 ( .ip1(n21179), .ip2(n22364), .ip3(n21120), .ip4(
        n20345), .op(n20349) );
  inv_1 U23242 ( .ip(n20346), .op(n20347) );
  nor2_1 U23243 ( .ip1(n22254), .ip2(n20347), .op(n20348) );
  nor2_1 U23244 ( .ip1(n20349), .ip2(n20348), .op(\pipeline/csr/N1943 ) );
  inv_1 U23245 ( .ip(n20350), .op(n20351) );
  nor2_1 U23246 ( .ip1(\pipeline/csr/mtime_full [6]), .ip2(n20351), .op(n20354) );
  nor3_1 U23247 ( .ip1(n21193), .ip2(n20353), .ip3(n20354), .op(n20352) );
  not_ab_or_c_or_d U23248 ( .ip1(n21195), .ip2(n22364), .ip3(n21217), .ip4(
        n20352), .op(n20357) );
  nor2_1 U23249 ( .ip1(n20354), .ip2(n20353), .op(n20355) );
  nor2_1 U23250 ( .ip1(n21198), .ip2(n20355), .op(n20356) );
  nor2_1 U23251 ( .ip1(n20357), .ip2(n20356), .op(\pipeline/csr/N2087 ) );
  nand2_1 U23252 ( .ip1(n22013), .ip2(\pipeline/csr/mscratch [6]), .op(n20359)
         );
  nand2_1 U23253 ( .ip1(n22014), .ip2(n22364), .op(n20358) );
  nand2_1 U23254 ( .ip1(n20359), .ip2(n20358), .op(n9922) );
  nand2_1 U23255 ( .ip1(n22372), .ip2(\pipeline/csr/from_host [6]), .op(n20361) );
  nand2_1 U23256 ( .ip1(n22373), .ip2(n22364), .op(n20360) );
  nand2_1 U23257 ( .ip1(n20361), .ip2(n20360), .op(n9954) );
  nand2_1 U23258 ( .ip1(n22378), .ip2(n22364), .op(n20363) );
  nand2_1 U23259 ( .ip1(n22376), .ip2(\pipeline/csr/to_host [6]), .op(n20362)
         );
  nand2_1 U23260 ( .ip1(n20363), .ip2(n20362), .op(n8766) );
  or2_1 U23261 ( .ip1(\pipeline/csr/cycle_full [6]), .ip2(n21077), .op(n20364)
         );
  nand2_1 U23262 ( .ip1(n20365), .ip2(n20364), .op(n20366) );
  or2_1 U23263 ( .ip1(n21145), .ip2(n20366), .op(n20368) );
  nand2_1 U23264 ( .ip1(n22021), .ip2(n22364), .op(n20367) );
  nand2_1 U23265 ( .ip1(n20368), .ip2(n20367), .op(\pipeline/csr/N1879 ) );
  nor2_1 U23266 ( .ip1(n20990), .ip2(n20370), .op(n20373) );
  not_ab_or_c_or_d U23267 ( .ip1(n20371), .ip2(n20370), .ip3(n21005), .ip4(
        n20369), .op(n20372) );
  ab_or_c_or_d U23268 ( .ip1(n21019), .ip2(n22364), .ip3(n20373), .ip4(n20372), 
        .op(n10132) );
  nand2_1 U23269 ( .ip1(n22314), .ip2(n22364), .op(n20377) );
  or2_1 U23270 ( .ip1(\pipeline/csr/cycle_full [38]), .ip2(n21068), .op(n20374) );
  nand3_1 U23271 ( .ip1(n20375), .ip2(n20374), .ip3(n22316), .op(n20376) );
  nand2_1 U23272 ( .ip1(n20377), .ip2(n20376), .op(\pipeline/csr/N1911 ) );
  inv_1 U23273 ( .ip(n20378), .op(n20379) );
  mux2_1 U23274 ( .ip1(\pipeline/csr_rdata_WB [6]), .ip2(n20379), .s(n20389), 
        .op(n8800) );
  xor2_1 U23275 ( .ip1(n20381), .ip2(n20380), .op(n20382) );
  nand2_1 U23276 ( .ip1(n21649), .ip2(n20382), .op(n20388) );
  nor2_1 U23277 ( .ip1(\pipeline/md/b [7]), .ip2(n20384), .op(n20383) );
  not_ab_or_c_or_d U23278 ( .ip1(\pipeline/md/b [7]), .ip2(n20384), .ip3(
        n21884), .ip4(n20383), .op(n20385) );
  xor2_1 U23279 ( .ip1(\pipeline/md/a [7]), .ip2(n20385), .op(n20386) );
  nand2_1 U23280 ( .ip1(n20386), .ip2(n21643), .op(n20387) );
  nand2_1 U23281 ( .ip1(n20388), .ip2(n20387), .op(n8373) );
  mux2_1 U23282 ( .ip1(\pipeline/csr_rdata_WB [7]), .ip2(n20390), .s(n20389), 
        .op(n8799) );
  xor2_1 U23283 ( .ip1(n20392), .ip2(n20391), .op(n20393) );
  nand2_1 U23284 ( .ip1(n21649), .ip2(n20393), .op(n20398) );
  xor2_1 U23285 ( .ip1(\pipeline/md/b [12]), .ip2(n20403), .op(n20394) );
  nor2_1 U23286 ( .ip1(n21884), .ip2(n20394), .op(n20395) );
  xor2_1 U23287 ( .ip1(\pipeline/md/a [12]), .ip2(n20395), .op(n20396) );
  nand2_1 U23288 ( .ip1(n20396), .ip2(n21643), .op(n20397) );
  nand2_1 U23289 ( .ip1(n20398), .ip2(n20397), .op(n8411) );
  xor2_1 U23290 ( .ip1(n20400), .ip2(n20399), .op(n20401) );
  nand2_1 U23291 ( .ip1(n21649), .ip2(n20401), .op(n20409) );
  and2_1 U23292 ( .ip1(n20403), .ip2(n20402), .op(n20413) );
  nor2_1 U23293 ( .ip1(n20413), .ip2(n20412), .op(n20405) );
  nor2_1 U23294 ( .ip1(\pipeline/md/b [13]), .ip2(n20405), .op(n20404) );
  not_ab_or_c_or_d U23295 ( .ip1(\pipeline/md/b [13]), .ip2(n20405), .ip3(
        n21884), .ip4(n20404), .op(n20406) );
  xor2_1 U23296 ( .ip1(\pipeline/md/a [13]), .ip2(n20406), .op(n20407) );
  nand2_1 U23297 ( .ip1(n20407), .ip2(n21643), .op(n20408) );
  nand2_1 U23298 ( .ip1(n20409), .ip2(n20408), .op(n8406) );
  xor2_1 U23299 ( .ip1(n20424), .ip2(n20423), .op(n20410) );
  nand2_1 U23300 ( .ip1(n21649), .ip2(n20410), .op(n20422) );
  or3_1 U23301 ( .ip1(n20413), .ip2(n20412), .ip3(n20411), .op(n20415) );
  nand2_1 U23302 ( .ip1(n20415), .ip2(n20414), .op(n20416) );
  xor2_1 U23303 ( .ip1(n20417), .ip2(n20416), .op(n20418) );
  nor2_1 U23304 ( .ip1(n21947), .ip2(n20418), .op(n20419) );
  xor2_1 U23305 ( .ip1(\pipeline/md/a [14]), .ip2(n20419), .op(n20420) );
  nand2_1 U23306 ( .ip1(n20420), .ip2(n21643), .op(n20421) );
  nand2_1 U23307 ( .ip1(n20422), .ip2(n20421), .op(n8389) );
  nand2_1 U23308 ( .ip1(n20424), .ip2(n20423), .op(n20425) );
  nand2_1 U23309 ( .ip1(n20426), .ip2(n20425), .op(n20427) );
  nand2_1 U23310 ( .ip1(n21649), .ip2(n20427), .op(n20428) );
  nand2_1 U23311 ( .ip1(n20649), .ip2(n20428), .op(n20429) );
  nand2_1 U23312 ( .ip1(n20430), .ip2(n20429), .op(n20439) );
  inv_1 U23313 ( .ip(n20431), .op(n20432) );
  nor2_1 U23314 ( .ip1(n20433), .ip2(n20432), .op(n20434) );
  xor2_1 U23315 ( .ip1(\pipeline/md/b [15]), .ip2(n20434), .op(n20435) );
  nor2_1 U23316 ( .ip1(n21947), .ip2(n20435), .op(n20436) );
  xor2_1 U23317 ( .ip1(\pipeline/md/a [15]), .ip2(n20436), .op(n20437) );
  nand2_1 U23318 ( .ip1(n20437), .ip2(n21643), .op(n20438) );
  nand2_1 U23319 ( .ip1(n20439), .ip2(n20438), .op(n8382) );
  nor2_1 U23320 ( .ip1(n20440), .ip2(n20483), .op(n20441) );
  xor2_1 U23321 ( .ip1(n20441), .ip2(n15597), .op(n20442) );
  nand2_1 U23322 ( .ip1(n21649), .ip2(n20442), .op(n20448) );
  xor2_1 U23323 ( .ip1(\pipeline/md/b [18]), .ip2(n20443), .op(n20444) );
  nor2_1 U23324 ( .ip1(n21947), .ip2(n20444), .op(n20445) );
  xor2_1 U23325 ( .ip1(\pipeline/md/a [18]), .ip2(n20445), .op(n20446) );
  nand2_1 U23326 ( .ip1(n20446), .ip2(n21643), .op(n20447) );
  nand2_1 U23327 ( .ip1(n20448), .ip2(n20447), .op(n8396) );
  nor4_1 U23328 ( .ip1(\pipeline/md_resp_result [21]), .ip2(n20463), .ip3(
        n20462), .ip4(n22755), .op(n20460) );
  nand2_1 U23329 ( .ip1(\pipeline/md/negate_output ), .ip2(n20449), .op(n20451) );
  nor2_1 U23330 ( .ip1(n20452), .ip2(n20451), .op(n20450) );
  not_ab_or_c_or_d U23331 ( .ip1(n20452), .ip2(n20451), .ip3(n21960), .ip4(
        n20450), .op(n20458) );
  nor3_1 U23332 ( .ip1(\pipeline/md/result [53]), .ip2(n20453), .ip3(n21966), 
        .op(n20456) );
  inv_1 U23333 ( .ip(n20453), .op(n20454) );
  not_ab_or_c_or_d U23334 ( .ip1(\pipeline/md/negate_output ), .ip2(n20454), 
        .ip3(n22679), .ip4(n21967), .op(n20455) );
  nor3_1 U23335 ( .ip1(n21972), .ip2(n20456), .ip3(n20455), .op(n20457) );
  nor2_1 U23336 ( .ip1(n20458), .ip2(n20457), .op(n20459) );
  not_ab_or_c_or_d U23337 ( .ip1(n20680), .ip2(n20461), .ip3(n20460), .ip4(
        n20459), .op(n20468) );
  or2_1 U23338 ( .ip1(n20463), .ip2(n20462), .op(n20464) );
  nand2_1 U23339 ( .ip1(n21440), .ip2(n20464), .op(n20465) );
  nand2_1 U23340 ( .ip1(n22738), .ip2(n20465), .op(n20466) );
  nand2_1 U23341 ( .ip1(\pipeline/md_resp_result [21]), .ip2(n20466), .op(
        n20467) );
  nand2_1 U23342 ( .ip1(n20468), .ip2(n20467), .op(n8613) );
  mux2_1 U23343 ( .ip1(\pipeline/csr_rdata_WB [21]), .ip2(n20469), .s(n17429), 
        .op(n8785) );
  nand2_1 U23344 ( .ip1(n21995), .ip2(imem_haddr[22]), .op(n20471) );
  nand2_1 U23345 ( .ip1(\pipeline/PC_IF [22]), .ip2(n21996), .op(n20470) );
  nand2_1 U23346 ( .ip1(n20471), .ip2(n20470), .op(n8446) );
  nand2_1 U23347 ( .ip1(\pipeline/PC_IF [22]), .ip2(n22048), .op(n20473) );
  nand2_1 U23348 ( .ip1(\pipeline/PC_DX [22]), .ip2(n21999), .op(n20472) );
  nand2_1 U23349 ( .ip1(n20473), .ip2(n20472), .op(n8445) );
  mux2_1 U23350 ( .ip1(dmem_haddr[5]), .ip2(\pipeline/alu_out_WB [5]), .s(
        n19505), .op(n8727) );
  nand2_1 U23351 ( .ip1(n21624), .ip2(n20474), .op(n20475) );
  xor2_1 U23352 ( .ip1(n20476), .ip2(n20475), .op(n20477) );
  nor2_1 U23353 ( .ip1(n20477), .ip2(n21499), .op(n20482) );
  xor2_1 U23354 ( .ip1(\pipeline/md/a [5]), .ip2(\pipeline/md/b [5]), .op(
        n20478) );
  xor2_1 U23355 ( .ip1(n20479), .ip2(n20478), .op(n20480) );
  nor2_1 U23356 ( .ip1(n20480), .ip2(n21730), .op(n20481) );
  ab_or_c_or_d U23357 ( .ip1(\pipeline/md/a [5]), .ip2(n21947), .ip3(n20482), 
        .ip4(n20481), .op(n8378) );
  nor2_1 U23358 ( .ip1(n20484), .ip2(n20483), .op(n20486) );
  xor2_1 U23359 ( .ip1(n20486), .ip2(n20485), .op(n20487) );
  nand2_1 U23360 ( .ip1(n21649), .ip2(n20487), .op(n20493) );
  xor2_1 U23361 ( .ip1(\pipeline/md/b [6]), .ip2(n20488), .op(n20489) );
  nor2_1 U23362 ( .ip1(n21947), .ip2(n20489), .op(n20490) );
  xor2_1 U23363 ( .ip1(\pipeline/md/a [6]), .ip2(n20490), .op(n20491) );
  nand2_1 U23364 ( .ip1(n20491), .ip2(n21643), .op(n20492) );
  nand2_1 U23365 ( .ip1(n20493), .ip2(n20492), .op(n8366) );
  xor2_1 U23366 ( .ip1(n20507), .ip2(n20506), .op(n20494) );
  nand2_1 U23367 ( .ip1(n21649), .ip2(n20494), .op(n20505) );
  nand2_1 U23368 ( .ip1(n20496), .ip2(n20495), .op(n20498) );
  nand2_1 U23369 ( .ip1(n20498), .ip2(n20497), .op(n20499) );
  xor2_1 U23370 ( .ip1(n20500), .ip2(n20499), .op(n20501) );
  nor2_1 U23371 ( .ip1(n21947), .ip2(n20501), .op(n20502) );
  xor2_1 U23372 ( .ip1(\pipeline/md/a [9]), .ip2(n20502), .op(n20503) );
  nand2_1 U23373 ( .ip1(n20503), .ip2(n21643), .op(n20504) );
  nand2_1 U23374 ( .ip1(n20505), .ip2(n20504), .op(n8375) );
  inv_1 U23375 ( .ip(n20522), .op(n20512) );
  nand2_1 U23376 ( .ip1(n20507), .ip2(n20506), .op(n20508) );
  nand2_1 U23377 ( .ip1(n14601), .ip2(n20508), .op(n20509) );
  nand2_1 U23378 ( .ip1(n21649), .ip2(n20509), .op(n20510) );
  nand2_1 U23379 ( .ip1(n20649), .ip2(n20510), .op(n20511) );
  nand2_1 U23380 ( .ip1(n20512), .ip2(n20511), .op(n20520) );
  nor2_1 U23381 ( .ip1(n20514), .ip2(n20513), .op(n20527) );
  xor2_1 U23382 ( .ip1(n20527), .ip2(n20515), .op(n20516) );
  nor2_1 U23383 ( .ip1(n21947), .ip2(n20516), .op(n20517) );
  xor2_1 U23384 ( .ip1(\pipeline/md/a [10]), .ip2(n20517), .op(n20518) );
  nand2_1 U23385 ( .ip1(n20518), .ip2(n21643), .op(n20519) );
  nand2_1 U23386 ( .ip1(n20520), .ip2(n20519), .op(n8414) );
  nand2_1 U23387 ( .ip1(n21649), .ip2(n20522), .op(n20521) );
  nand2_1 U23388 ( .ip1(n20649), .ip2(n20521), .op(n20525) );
  nor2_1 U23389 ( .ip1(n20522), .ip2(n20647), .op(n20524) );
  mux2_1 U23390 ( .ip1(n20525), .ip2(n20524), .s(n20523), .op(n20536) );
  nor2_1 U23391 ( .ip1(n20527), .ip2(n20526), .op(n20530) );
  inv_1 U23392 ( .ip(n20528), .op(n20529) );
  nor2_1 U23393 ( .ip1(n20530), .ip2(n20529), .op(n20531) );
  xor2_1 U23394 ( .ip1(\pipeline/md/b [11]), .ip2(n20531), .op(n20532) );
  nand2_1 U23395 ( .ip1(n20532), .ip2(n14770), .op(n20533) );
  xor2_1 U23396 ( .ip1(\pipeline/md/a [11]), .ip2(n20533), .op(n20534) );
  nor2_1 U23397 ( .ip1(n21866), .ip2(n20534), .op(n20535) );
  or2_1 U23398 ( .ip1(n20536), .ip2(n20535), .op(n8420) );
  nor3_1 U23399 ( .ip1(n20537), .ip2(n20544), .ip3(n21957), .op(n20542) );
  nor2_1 U23400 ( .ip1(n20538), .ip2(n21659), .op(n20540) );
  nor2_1 U23401 ( .ip1(\pipeline/md/result [51]), .ip2(n20540), .op(n20539) );
  not_ab_or_c_or_d U23402 ( .ip1(\pipeline/md/result [51]), .ip2(n20540), 
        .ip3(n21662), .ip4(n20539), .op(n20541) );
  or2_1 U23403 ( .ip1(n20542), .ip2(n20541), .op(n20551) );
  nand2_1 U23404 ( .ip1(n21972), .ip2(n20543), .op(n20548) );
  nand2_1 U23405 ( .ip1(n20552), .ip2(n20669), .op(n20547) );
  inv_1 U23406 ( .ip(n20544), .op(n20545) );
  not_ab_or_c_or_d U23407 ( .ip1(n20548), .ip2(n20547), .ip3(n20546), .ip4(
        n20545), .op(n20550) );
  nor4_1 U23408 ( .ip1(\pipeline/md_resp_result [19]), .ip2(n20556), .ip3(
        n20555), .ip4(n22755), .op(n20549) );
  not_ab_or_c_or_d U23409 ( .ip1(n20552), .ip2(n20551), .ip3(n20550), .ip4(
        n20549), .op(n20562) );
  nand2_1 U23410 ( .ip1(n20554), .ip2(n20553), .op(n20561) );
  or2_1 U23411 ( .ip1(n20556), .ip2(n20555), .op(n20557) );
  nand2_1 U23412 ( .ip1(n21440), .ip2(n20557), .op(n20558) );
  nand2_1 U23413 ( .ip1(n22738), .ip2(n20558), .op(n20559) );
  nand2_1 U23414 ( .ip1(\pipeline/md_resp_result [19]), .ip2(n20559), .op(
        n20560) );
  nand3_1 U23415 ( .ip1(n20562), .ip2(n20561), .ip3(n20560), .op(n8615) );
  mux2_1 U23416 ( .ip1(\pipeline/csr_rdata_WB [19]), .ip2(n20563), .s(n17777), 
        .op(n8787) );
  nand2_1 U23417 ( .ip1(n20565), .ip2(n20564), .op(n20566) );
  xor2_1 U23418 ( .ip1(\pipeline/md/b [19]), .ip2(n20566), .op(n20567) );
  nor2_1 U23419 ( .ip1(n21947), .ip2(n20567), .op(n20568) );
  xor2_1 U23420 ( .ip1(\pipeline/md/a [19]), .ip2(n20568), .op(n20569) );
  nand2_1 U23421 ( .ip1(n20569), .ip2(n21643), .op(n20574) );
  xor2_1 U23422 ( .ip1(n20571), .ip2(n20570), .op(n20572) );
  nand2_1 U23423 ( .ip1(n21649), .ip2(n20572), .op(n20573) );
  nand2_1 U23424 ( .ip1(n20574), .ip2(n20573), .op(n8391) );
  xor2_1 U23425 ( .ip1(n20584), .ip2(n20583), .op(n20575) );
  nand2_1 U23426 ( .ip1(n21649), .ip2(n20575), .op(n20582) );
  xor2_1 U23427 ( .ip1(n20577), .ip2(n20576), .op(n20578) );
  nor2_1 U23428 ( .ip1(n21884), .ip2(n20578), .op(n20579) );
  xor2_1 U23429 ( .ip1(\pipeline/md/a [20]), .ip2(n20579), .op(n20580) );
  nand2_1 U23430 ( .ip1(n20580), .ip2(n21643), .op(n20581) );
  nand2_1 U23431 ( .ip1(n20582), .ip2(n20581), .op(n8410) );
  nand2_1 U23432 ( .ip1(n20584), .ip2(n20583), .op(n20585) );
  nand2_1 U23433 ( .ip1(n20586), .ip2(n20585), .op(n20587) );
  nand2_1 U23434 ( .ip1(n21649), .ip2(n20587), .op(n20588) );
  nand2_1 U23435 ( .ip1(n20649), .ip2(n20588), .op(n20589) );
  nand2_1 U23436 ( .ip1(n20598), .ip2(n20589), .op(n20596) );
  xor2_1 U23437 ( .ip1(n20591), .ip2(n20590), .op(n20592) );
  nor2_1 U23438 ( .ip1(n21947), .ip2(n20592), .op(n20593) );
  xor2_1 U23439 ( .ip1(\pipeline/md/a [21]), .ip2(n20593), .op(n20594) );
  nand2_1 U23440 ( .ip1(n20594), .ip2(n21643), .op(n20595) );
  nand2_1 U23441 ( .ip1(n20596), .ip2(n20595), .op(n8404) );
  nor2_1 U23442 ( .ip1(n21499), .ip2(n20598), .op(n20597) );
  nor2_1 U23443 ( .ip1(n20633), .ip2(n20597), .op(n20601) );
  nand2_1 U23444 ( .ip1(n20634), .ip2(n20598), .op(n20600) );
  mux2_1 U23445 ( .ip1(n20601), .ip2(n20600), .s(n20599), .op(n20608) );
  xor2_1 U23446 ( .ip1(n20603), .ip2(n20602), .op(n20604) );
  nor2_1 U23447 ( .ip1(n21884), .ip2(n20604), .op(n20605) );
  xor2_1 U23448 ( .ip1(\pipeline/md/a [22]), .ip2(n20605), .op(n20606) );
  nand2_1 U23449 ( .ip1(n20606), .ip2(n21643), .op(n20607) );
  nand2_1 U23450 ( .ip1(n20608), .ip2(n20607), .op(n8409) );
  nor2_1 U23451 ( .ip1(n20647), .ip2(n20609), .op(n20613) );
  nand2_1 U23452 ( .ip1(n20609), .ip2(n21649), .op(n20610) );
  nand2_1 U23453 ( .ip1(n20610), .ip2(n20649), .op(n20612) );
  mux2_1 U23454 ( .ip1(n20613), .ip2(n20612), .s(n20611), .op(n20621) );
  nor2_1 U23455 ( .ip1(n20616), .ip2(n20615), .op(n20614) );
  not_ab_or_c_or_d U23456 ( .ip1(n20616), .ip2(n20615), .ip3(n21884), .ip4(
        n20614), .op(n20618) );
  xor2_1 U23457 ( .ip1(n20618), .ip2(n20617), .op(n20619) );
  nor2_1 U23458 ( .ip1(n21866), .ip2(n20619), .op(n20620) );
  or2_1 U23459 ( .ip1(n20621), .ip2(n20620), .op(n8424) );
  nor2_1 U23460 ( .ip1(n20647), .ip2(n20622), .op(n20625) );
  nand2_1 U23461 ( .ip1(n20622), .ip2(n21649), .op(n20623) );
  nand2_1 U23462 ( .ip1(n20623), .ip2(n20649), .op(n20624) );
  mux2_1 U23463 ( .ip1(n20625), .ip2(n20624), .s(n16333), .op(n20631) );
  xor2_1 U23464 ( .ip1(\pipeline/md/b [26]), .ip2(n20626), .op(n20627) );
  nand2_1 U23465 ( .ip1(n14770), .ip2(n20627), .op(n20628) );
  xor2_1 U23466 ( .ip1(\pipeline/md/a [26]), .ip2(n20628), .op(n20629) );
  nor2_1 U23467 ( .ip1(n21866), .ip2(n20629), .op(n20630) );
  or2_1 U23468 ( .ip1(n20631), .ip2(n20630), .op(n8412) );
  nor2_1 U23469 ( .ip1(n21499), .ip2(n20645), .op(n20632) );
  nor2_1 U23470 ( .ip1(n20633), .ip2(n20632), .op(n20637) );
  nand2_1 U23471 ( .ip1(n20634), .ip2(n20645), .op(n20636) );
  mux2_1 U23472 ( .ip1(n20637), .ip2(n20636), .s(n20635), .op(n20644) );
  nor2_1 U23473 ( .ip1(n20639), .ip2(n20638), .op(n20654) );
  xor2_1 U23474 ( .ip1(n20654), .ip2(\pipeline/md/b [28]), .op(n20640) );
  nor2_1 U23475 ( .ip1(n21884), .ip2(n20640), .op(n20641) );
  xor2_1 U23476 ( .ip1(\pipeline/md/a [28]), .ip2(n20641), .op(n20642) );
  nand2_1 U23477 ( .ip1(n20642), .ip2(n21643), .op(n20643) );
  nand2_1 U23478 ( .ip1(n20644), .ip2(n20643), .op(n8423) );
  nor2_1 U23479 ( .ip1(n20646), .ip2(n20645), .op(n21621) );
  nor2_1 U23480 ( .ip1(n20647), .ip2(n21621), .op(n20652) );
  nand2_1 U23481 ( .ip1(n21621), .ip2(n21649), .op(n20648) );
  nand2_1 U23482 ( .ip1(n20649), .ip2(n20648), .op(n20651) );
  mux2_1 U23483 ( .ip1(n20652), .ip2(n20651), .s(n20650), .op(n20662) );
  nor2_1 U23484 ( .ip1(n20654), .ip2(n20653), .op(n20656) );
  nor2_1 U23485 ( .ip1(n20656), .ip2(n20655), .op(n21628) );
  xor2_1 U23486 ( .ip1(n21628), .ip2(n20657), .op(n20658) );
  nand2_1 U23487 ( .ip1(n14770), .ip2(n20658), .op(n20659) );
  xor2_1 U23488 ( .ip1(\pipeline/md/a [29]), .ip2(n20659), .op(n20660) );
  nor2_1 U23489 ( .ip1(n21866), .ip2(n20660), .op(n20661) );
  or2_1 U23490 ( .ip1(n20662), .ip2(n20661), .op(n8415) );
  nor4_1 U23491 ( .ip1(\pipeline/md_resp_result [29]), .ip2(n20682), .ip3(
        n20681), .ip4(n22755), .op(n20679) );
  nor2_1 U23492 ( .ip1(n20666), .ip2(n21659), .op(n20663) );
  nor2_1 U23493 ( .ip1(n20664), .ip2(n20663), .op(n20671) );
  inv_1 U23494 ( .ip(n20664), .op(n20665) );
  nor2_1 U23495 ( .ip1(n20666), .ip2(n20665), .op(n20667) );
  nor2_1 U23496 ( .ip1(n21960), .ip2(n20667), .op(n20668) );
  nor2_1 U23497 ( .ip1(n20669), .ip2(n20668), .op(n20670) );
  nor2_1 U23498 ( .ip1(n20671), .ip2(n20670), .op(n20677) );
  nor3_1 U23499 ( .ip1(\pipeline/md/result [61]), .ip2(n20672), .ip3(n21966), 
        .op(n20675) );
  inv_1 U23500 ( .ip(n20672), .op(n20673) );
  not_ab_or_c_or_d U23501 ( .ip1(\pipeline/md/negate_output ), .ip2(n20673), 
        .ip3(n22743), .ip4(n21967), .op(n20674) );
  nor3_1 U23502 ( .ip1(n21972), .ip2(n20675), .ip3(n20674), .op(n20676) );
  nor2_1 U23503 ( .ip1(n20677), .ip2(n20676), .op(n20678) );
  not_ab_or_c_or_d U23504 ( .ip1(n20680), .ip2(n21672), .ip3(n20679), .ip4(
        n20678), .op(n20687) );
  or2_1 U23505 ( .ip1(n20682), .ip2(n20681), .op(n20683) );
  nand2_1 U23506 ( .ip1(n21440), .ip2(n20683), .op(n20684) );
  nand2_1 U23507 ( .ip1(n22738), .ip2(n20684), .op(n20685) );
  nand2_1 U23508 ( .ip1(\pipeline/md_resp_result [29]), .ip2(n20685), .op(
        n20686) );
  nand2_1 U23509 ( .ip1(n20687), .ip2(n20686), .op(n8605) );
  mux2_1 U23510 ( .ip1(\pipeline/csr_rdata_WB [29]), .ip2(n20688), .s(n19498), 
        .op(n8777) );
  nand2_1 U23511 ( .ip1(n20690), .ip2(n20689), .op(n20694) );
  nor2_1 U23512 ( .ip1(n20692), .ip2(n20691), .op(n20693) );
  xor2_1 U23513 ( .ip1(n20694), .ip2(n20693), .op(imem_haddr[11]) );
  nand2_1 U23514 ( .ip1(n21995), .ip2(imem_haddr[11]), .op(n20696) );
  nand2_1 U23515 ( .ip1(\pipeline/PC_IF [11]), .ip2(n21996), .op(n20695) );
  nand2_1 U23516 ( .ip1(n20696), .ip2(n20695), .op(n8468) );
  nand2_1 U23517 ( .ip1(\pipeline/PC_IF [11]), .ip2(n21988), .op(n20698) );
  nand2_1 U23518 ( .ip1(\pipeline/PC_DX [11]), .ip2(n21999), .op(n20697) );
  nand2_1 U23519 ( .ip1(n20698), .ip2(n20697), .op(n8467) );
  mux2_1 U23520 ( .ip1(\pipeline/PC_WB [11]), .ip2(\pipeline/PC_DX [11]), .s(
        n19498), .op(n8892) );
  nand2_1 U23521 ( .ip1(n20788), .ip2(n21043), .op(n20704) );
  and2_1 U23522 ( .ip1(n21174), .ip2(\pipeline/epc [12]), .op(n20702) );
  xor2_1 U23523 ( .ip1(\pipeline/PC_WB [12]), .ip2(n20699), .op(n20700) );
  nor2_1 U23524 ( .ip1(n21171), .ip2(n20700), .op(n20701) );
  nor2_1 U23525 ( .ip1(n20702), .ip2(n20701), .op(n20703) );
  nand2_1 U23526 ( .ip1(n20704), .ip2(n20703), .op(n8859) );
  nand2_1 U23527 ( .ip1(n21032), .ip2(n20788), .op(n20707) );
  nand2_1 U23528 ( .ip1(\pipeline/csr/mtvec [12]), .ip2(n20705), .op(n20706)
         );
  nand2_1 U23529 ( .ip1(n20707), .ip2(n20706), .op(n9980) );
  nand2_1 U23530 ( .ip1(n20709), .ip2(n20708), .op(n20722) );
  inv_1 U23531 ( .ip(n20710), .op(n20714) );
  nor2_1 U23532 ( .ip1(n20712), .ip2(n20711), .op(n20713) );
  nor2_1 U23533 ( .ip1(n20714), .ip2(n20713), .op(n20720) );
  nand2_1 U23534 ( .ip1(n20716), .ip2(n20715), .op(n20718) );
  or2_1 U23535 ( .ip1(n20718), .ip2(n20717), .op(n20719) );
  nand2_1 U23536 ( .ip1(n20720), .ip2(n20719), .op(n20721) );
  xnor2_1 U23537 ( .ip1(n20722), .ip2(n20721), .op(n20744) );
  nor2_1 U23538 ( .ip1(n20724), .ip2(n20723), .op(n20743) );
  or2_1 U23539 ( .ip1(n20726), .ip2(n20725), .op(n20741) );
  nand2_1 U23540 ( .ip1(n10189), .ip2(n20727), .op(n20732) );
  and3_1 U23541 ( .ip1(n13627), .ip2(n20904), .ip3(n20728), .op(n20731) );
  nor2_1 U23542 ( .ip1(n21555), .ip2(n20729), .op(n20730) );
  not_ab_or_c_or_d U23543 ( .ip1(n21557), .ip2(n20732), .ip3(n20731), .ip4(
        n20730), .op(n20740) );
  nand2_1 U23544 ( .ip1(n20733), .ip2(n21544), .op(n20734) );
  mux2_1 U23545 ( .ip1(n20735), .ip2(n20734), .s(n19427), .op(n20739) );
  nand2_1 U23546 ( .ip1(n20737), .ip2(n20736), .op(n20738) );
  ab_or_c_or_d U23547 ( .ip1(n20744), .ip2(n21577), .ip3(n20743), .ip4(n20742), 
        .op(dmem_haddr[12]) );
  mux2_1 U23548 ( .ip1(dmem_haddr[12]), .ip2(\pipeline/alu_out_WB [12]), .s(
        n21582), .op(n8720) );
  inv_1 U23549 ( .ip(\pipeline/csr/time_full [44]), .op(n20746) );
  nor2_1 U23550 ( .ip1(n20747), .ip2(n20746), .op(n20745) );
  not_ab_or_c_or_d U23551 ( .ip1(n20747), .ip2(n20746), .ip3(n22282), .ip4(
        n20745), .op(n20751) );
  inv_1 U23552 ( .ip(n20788), .op(n22161) );
  nor2_1 U23553 ( .ip1(n22161), .ip2(n20748), .op(n20749) );
  nor2_1 U23554 ( .ip1(n20749), .ip2(n22284), .op(n20750) );
  nor2_1 U23555 ( .ip1(n20751), .ip2(n20750), .op(\pipeline/csr/N1981 ) );
  or2_1 U23556 ( .ip1(\pipeline/csr/time_full [12]), .ip2(n20752), .op(n20753)
         );
  nand2_1 U23557 ( .ip1(n20754), .ip2(n20753), .op(n20755) );
  or2_1 U23558 ( .ip1(n22002), .ip2(n20755), .op(n20757) );
  nand2_1 U23559 ( .ip1(n22005), .ip2(n20788), .op(n20756) );
  nand2_1 U23560 ( .ip1(n20757), .ip2(n20756), .op(\pipeline/csr/N1949 ) );
  inv_1 U23561 ( .ip(n20758), .op(n20759) );
  nor2_1 U23562 ( .ip1(\pipeline/csr/mtime_full [12]), .ip2(n20759), .op(
        n20762) );
  nor3_1 U23563 ( .ip1(n21193), .ip2(n20762), .ip3(n20761), .op(n20760) );
  not_ab_or_c_or_d U23564 ( .ip1(n21195), .ip2(n20788), .ip3(n21120), .ip4(
        n20760), .op(n20765) );
  nor2_1 U23565 ( .ip1(n20762), .ip2(n20761), .op(n20763) );
  nor2_1 U23566 ( .ip1(n22254), .ip2(n20763), .op(n20764) );
  nor2_1 U23567 ( .ip1(n20765), .ip2(n20764), .op(\pipeline/csr/N2093 ) );
  nand2_1 U23568 ( .ip1(\pipeline/csr/mscratch [12]), .ip2(n22013), .op(n20767) );
  nand2_1 U23569 ( .ip1(n22014), .ip2(n20788), .op(n20766) );
  nand2_1 U23570 ( .ip1(n20767), .ip2(n20766), .op(n9916) );
  nand2_1 U23571 ( .ip1(\pipeline/csr/from_host [12]), .ip2(n22372), .op(
        n20769) );
  nand2_1 U23572 ( .ip1(n22373), .ip2(n20788), .op(n20768) );
  nand2_1 U23573 ( .ip1(n20769), .ip2(n20768), .op(n9948) );
  nand2_1 U23574 ( .ip1(n22378), .ip2(n20788), .op(n20771) );
  nand2_1 U23575 ( .ip1(\pipeline/csr/to_host [12]), .ip2(n22376), .op(n20770)
         );
  nand2_1 U23576 ( .ip1(n20771), .ip2(n20770), .op(n8760) );
  or2_1 U23577 ( .ip1(\pipeline/csr/cycle_full [12]), .ip2(n20772), .op(n20773) );
  nand2_1 U23578 ( .ip1(n20774), .ip2(n20773), .op(n20775) );
  or2_1 U23579 ( .ip1(n21145), .ip2(n20775), .op(n20777) );
  nand2_1 U23580 ( .ip1(n22021), .ip2(n20788), .op(n20776) );
  nand2_1 U23581 ( .ip1(n20777), .ip2(n20776), .op(\pipeline/csr/N1885 ) );
  nand2_1 U23582 ( .ip1(\pipeline/csr/mtimecmp [12]), .ip2(n22363), .op(n20779) );
  nand2_1 U23583 ( .ip1(n22365), .ip2(n20788), .op(n20778) );
  nand2_1 U23584 ( .ip1(n20779), .ip2(n20778), .op(n10010) );
  nand2_1 U23585 ( .ip1(n21019), .ip2(n20788), .op(n20785) );
  nand2_1 U23586 ( .ip1(\pipeline/csr/instret_full [12]), .ip2(n21016), .op(
        n20784) );
  mux2_1 U23587 ( .ip1(\pipeline/csr/instret_full [12]), .ip2(n20781), .s(
        n20780), .op(n20782) );
  or2_1 U23588 ( .ip1(n20782), .ip2(n21005), .op(n20783) );
  nand3_1 U23589 ( .ip1(n20785), .ip2(n20784), .ip3(n20783), .op(n10126) );
  nand2_1 U23590 ( .ip1(\pipeline/csr/mie [12]), .ip2(n22356), .op(n20787) );
  nand2_1 U23591 ( .ip1(n22357), .ip2(n20788), .op(n20786) );
  nand2_1 U23592 ( .ip1(n20787), .ip2(n20786), .op(n10048) );
  nand2_1 U23593 ( .ip1(n22314), .ip2(n20788), .op(n20793) );
  or2_1 U23594 ( .ip1(\pipeline/csr/cycle_full [44]), .ip2(n20789), .op(n20790) );
  nand3_1 U23595 ( .ip1(n20791), .ip2(n20790), .ip3(n22316), .op(n20792) );
  nand2_1 U23596 ( .ip1(n20793), .ip2(n20792), .op(\pipeline/csr/N1917 ) );
  inv_1 U23597 ( .ip(n20794), .op(n20795) );
  mux2_1 U23598 ( .ip1(\pipeline/csr_rdata_WB [12]), .ip2(n20795), .s(n17429), 
        .op(n8794) );
  xnor2_1 U23599 ( .ip1(n20797), .ip2(n20796), .op(imem_haddr[12]) );
  nand2_1 U23600 ( .ip1(n21995), .ip2(imem_haddr[12]), .op(n20799) );
  nand2_1 U23601 ( .ip1(\pipeline/PC_IF [12]), .ip2(n21996), .op(n20798) );
  nand2_1 U23602 ( .ip1(n20799), .ip2(n20798), .op(n8466) );
  nand2_1 U23603 ( .ip1(\pipeline/PC_IF [12]), .ip2(n22048), .op(n20801) );
  nand2_1 U23604 ( .ip1(\pipeline/PC_DX [12]), .ip2(n21999), .op(n20800) );
  nand2_1 U23605 ( .ip1(n20801), .ip2(n20800), .op(n8465) );
  mux2_1 U23606 ( .ip1(dmem_haddr[4]), .ip2(\pipeline/alu_out_WB [4]), .s(
        n21582), .op(n8728) );
  nand2_1 U23607 ( .ip1(n22282), .ip2(n22360), .op(n20804) );
  or2_1 U23608 ( .ip1(\pipeline/csr/time_full [36]), .ip2(n22269), .op(n20802)
         );
  nand3_1 U23609 ( .ip1(n21052), .ip2(n20802), .ip3(n22284), .op(n20803) );
  nand2_1 U23610 ( .ip1(n20804), .ip2(n20803), .op(\pipeline/csr/N1973 ) );
  inv_1 U23611 ( .ip(n21223), .op(n22268) );
  nor2_1 U23612 ( .ip1(n22268), .ip2(n21110), .op(n20808) );
  inv_1 U23613 ( .ip(n20811), .op(n20806) );
  nor2_1 U23614 ( .ip1(\pipeline/csr/instret_full [35]), .ip2(n21112), .op(
        n20805) );
  nor3_1 U23615 ( .ip1(n21111), .ip2(n20806), .ip3(n20805), .op(n20807) );
  ab_or_c_or_d U23616 ( .ip1(n21117), .ip2(\pipeline/csr/instret_full [35]), 
        .ip3(n20808), .ip4(n20807), .op(n10103) );
  nor2_1 U23617 ( .ip1(n19134), .ip2(n20810), .op(n20813) );
  not_ab_or_c_or_d U23618 ( .ip1(n20811), .ip2(n20810), .ip3(n21111), .ip4(
        n20809), .op(n20812) );
  ab_or_c_or_d U23619 ( .ip1(n20844), .ip2(n22360), .ip3(n20813), .ip4(n20812), 
        .op(n10102) );
  or2_1 U23620 ( .ip1(\pipeline/csr/time_full [4]), .ip2(n21180), .op(n20814)
         );
  nand2_1 U23621 ( .ip1(n21055), .ip2(n20814), .op(n20816) );
  nor2_1 U23622 ( .ip1(n21177), .ip2(n20816), .op(n20815) );
  not_ab_or_c_or_d U23623 ( .ip1(n21179), .ip2(n22360), .ip3(n21120), .ip4(
        n20815), .op(n20819) );
  inv_1 U23624 ( .ip(n20816), .op(n20817) );
  nor2_1 U23625 ( .ip1(n21198), .ip2(n20817), .op(n20818) );
  nor2_1 U23626 ( .ip1(n20819), .ip2(n20818), .op(\pipeline/csr/N1941 ) );
  inv_1 U23627 ( .ip(n20820), .op(n20821) );
  nor2_1 U23628 ( .ip1(\pipeline/csr/mtime_full [4]), .ip2(n20821), .op(n20823) );
  nor3_1 U23629 ( .ip1(n21193), .ip2(n21063), .ip3(n20823), .op(n20822) );
  not_ab_or_c_or_d U23630 ( .ip1(n21195), .ip2(n22360), .ip3(n21217), .ip4(
        n20822), .op(n20826) );
  nor2_1 U23631 ( .ip1(n20823), .ip2(n21063), .op(n20824) );
  nor2_1 U23632 ( .ip1(n22254), .ip2(n20824), .op(n20825) );
  nor2_1 U23633 ( .ip1(n20826), .ip2(n20825), .op(\pipeline/csr/N2085 ) );
  nand2_1 U23634 ( .ip1(n22013), .ip2(\pipeline/csr/mscratch [4]), .op(n20828)
         );
  nand2_1 U23635 ( .ip1(n22014), .ip2(n22360), .op(n20827) );
  nand2_1 U23636 ( .ip1(n20828), .ip2(n20827), .op(n9924) );
  nand2_1 U23637 ( .ip1(n22372), .ip2(\pipeline/csr/from_host [4]), .op(n20830) );
  nand2_1 U23638 ( .ip1(n22373), .ip2(n22360), .op(n20829) );
  nand2_1 U23639 ( .ip1(n20830), .ip2(n20829), .op(n9956) );
  nand2_1 U23640 ( .ip1(n22378), .ip2(n22360), .op(n20832) );
  nand2_1 U23641 ( .ip1(n22376), .ip2(\pipeline/csr/to_host [4]), .op(n20831)
         );
  nand2_1 U23642 ( .ip1(n20832), .ip2(n20831), .op(n8768) );
  or2_1 U23643 ( .ip1(\pipeline/csr/cycle_full [4]), .ip2(n21218), .op(n20833)
         );
  nand2_1 U23644 ( .ip1(n21073), .ip2(n20833), .op(n20834) );
  or2_1 U23645 ( .ip1(n21145), .ip2(n20834), .op(n20836) );
  nand2_1 U23646 ( .ip1(n22021), .ip2(n22360), .op(n20835) );
  nand2_1 U23647 ( .ip1(n20836), .ip2(n20835), .op(\pipeline/csr/N1877 ) );
  mux2_1 U23648 ( .ip1(\pipeline/PC_WB [0]), .ip2(\pipeline/PC_DX [0]), .s(
        n17777), .op(n8903) );
  nand2_1 U23649 ( .ip1(n22282), .ip2(n22377), .op(n20839) );
  or2_1 U23650 ( .ip1(\pipeline/csr/time_full [32]), .ip2(n20927), .op(n20837)
         );
  nand3_1 U23651 ( .ip1(n20837), .ip2(n22263), .ip3(n22284), .op(n20838) );
  nand2_1 U23652 ( .ip1(n20839), .ip2(n20838), .op(\pipeline/csr/N1969 ) );
  nor2_1 U23653 ( .ip1(n19134), .ip2(n20840), .op(n20843) );
  not_ab_or_c_or_d U23654 ( .ip1(n20841), .ip2(n20840), .ip3(n21111), .ip4(
        n21105), .op(n20842) );
  ab_or_c_or_d U23655 ( .ip1(n20844), .ip2(n22377), .ip3(n20843), .ip4(n20842), 
        .op(n10106) );
  or2_1 U23656 ( .ip1(n22002), .ip2(\pipeline/csr/time_full [0]), .op(n20846)
         );
  nand2_1 U23657 ( .ip1(n22005), .ip2(n22377), .op(n20845) );
  nand2_1 U23658 ( .ip1(n20846), .ip2(n20845), .op(\pipeline/csr/N1937 ) );
  mux2_1 U23659 ( .ip1(\pipeline/PC_WB [31]), .ip2(\pipeline/PC_DX [31]), .s(
        n20389), .op(n8872) );
  xor2_1 U23660 ( .ip1(\pipeline/PC_WB [31]), .ip2(n20847), .op(n20848) );
  nor2_1 U23661 ( .ip1(n21171), .ip2(n20848), .op(n20850) );
  nor2_1 U23662 ( .ip1(n22245), .ip2(n21168), .op(n20849) );
  ab_or_c_or_d U23663 ( .ip1(n21174), .ip2(\pipeline/epc [31]), .ip3(n20850), 
        .ip4(n20849), .op(n8840) );
  nor2_1 U23664 ( .ip1(n21029), .ip2(n20959), .op(n20854) );
  inv_1 U23665 ( .ip(\pipeline/csr/mtvec [31]), .op(n20851) );
  nor2_1 U23666 ( .ip1(n21089), .ip2(n20851), .op(n20852) );
  nor2_1 U23667 ( .ip1(n21032), .ip2(n20852), .op(n20853) );
  nor2_1 U23668 ( .ip1(n20854), .ip2(n20853), .op(n9961) );
  xor2_1 U23669 ( .ip1(n20903), .ip2(n20855), .op(n20857) );
  or2_1 U23670 ( .ip1(n20857), .ip2(n20856), .op(n20859) );
  nand2_1 U23671 ( .ip1(n20857), .ip2(n20856), .op(n20858) );
  nand2_1 U23672 ( .ip1(n20859), .ip2(n20858), .op(n20881) );
  nand2_1 U23673 ( .ip1(n20861), .ip2(n20860), .op(n20862) );
  nand2_1 U23674 ( .ip1(n20863), .ip2(n20862), .op(n20868) );
  nor2_1 U23675 ( .ip1(n20865), .ip2(n20864), .op(n20870) );
  and2_1 U23676 ( .ip1(n20866), .ip2(n20870), .op(n20867) );
  nor2_1 U23677 ( .ip1(n20868), .ip2(n20867), .op(n20873) );
  nand2_1 U23678 ( .ip1(n20870), .ip2(n20869), .op(n20875) );
  or2_1 U23679 ( .ip1(n20875), .ip2(n20871), .op(n20872) );
  nor2_1 U23680 ( .ip1(n20876), .ip2(n20875), .op(n20877) );
  nand2_1 U23681 ( .ip1(n20878), .ip2(n20877), .op(n20879) );
  nand2_1 U23682 ( .ip1(n20874), .ip2(n20879), .op(n20880) );
  xnor2_1 U23683 ( .ip1(n20881), .ip2(n20880), .op(n20919) );
  nor2_1 U23684 ( .ip1(n20883), .ip2(n20882), .op(n20918) );
  nor2_1 U23685 ( .ip1(n20885), .ip2(n20884), .op(n20889) );
  nor2_1 U23686 ( .ip1(n20887), .ip2(n20886), .op(n20888) );
  nor2_1 U23687 ( .ip1(n20889), .ip2(n20888), .op(n20901) );
  not_ab_or_c_or_d U23688 ( .ip1(n21536), .ip2(n20891), .ip3(n18918), .ip4(
        n20890), .op(n20895) );
  nand2_1 U23689 ( .ip1(n20892), .ip2(n17073), .op(n20893) );
  nand3_1 U23690 ( .ip1(n20895), .ip2(n20894), .ip3(n20893), .op(n20899) );
  nand2_1 U23691 ( .ip1(n20897), .ip2(n20896), .op(n20898) );
  nand4_1 U23692 ( .ip1(n20901), .ip2(n20900), .ip3(n20899), .ip4(n20898), 
        .op(n20916) );
  not_ab_or_c_or_d U23693 ( .ip1(n20904), .ip2(n20903), .ip3(n21557), .ip4(
        n20902), .op(n20906) );
  nor2_1 U23694 ( .ip1(n20906), .ip2(n20905), .op(n20909) );
  nor2_1 U23695 ( .ip1(n20907), .ip2(n10196), .op(n20908) );
  not_ab_or_c_or_d U23696 ( .ip1(n20911), .ip2(n20910), .ip3(n20909), .ip4(
        n20908), .op(n20915) );
  nand2_1 U23697 ( .ip1(n20913), .ip2(n20912), .op(n20914) );
  nand3_1 U23698 ( .ip1(n20916), .ip2(n20915), .ip3(n20914), .op(n20917) );
  ab_or_c_or_d U23699 ( .ip1(n20919), .ip2(n21577), .ip3(n20918), .ip4(n20917), 
        .op(dmem_haddr[31]) );
  mux2_1 U23700 ( .ip1(dmem_haddr[31]), .ip2(\pipeline/alu_out_WB [31]), .s(
        n21582), .op(n8701) );
  nor2_1 U23701 ( .ip1(n22245), .ip2(n21110), .op(n20922) );
  nor3_1 U23702 ( .ip1(n21111), .ip2(\pipeline/csr/instret_full [63]), .ip3(
        n20920), .op(n20921) );
  ab_or_c_or_d U23703 ( .ip1(\pipeline/csr/instret_full [63]), .ip2(n20923), 
        .ip3(n20922), .ip4(n20921), .op(n10075) );
  inv_1 U23704 ( .ip(n20924), .op(n20925) );
  nor2_1 U23705 ( .ip1(\pipeline/csr/time_full [31]), .ip2(n20925), .op(n20928) );
  nor3_1 U23706 ( .ip1(n21177), .ip2(n20927), .ip3(n20928), .op(n20926) );
  not_ab_or_c_or_d U23707 ( .ip1(n21179), .ip2(n20959), .ip3(n21217), .ip4(
        n20926), .op(n20931) );
  nor2_1 U23708 ( .ip1(n20928), .ip2(n20927), .op(n20929) );
  nor2_1 U23709 ( .ip1(n21198), .ip2(n20929), .op(n20930) );
  nor2_1 U23710 ( .ip1(n20931), .ip2(n20930), .op(\pipeline/csr/N1968 ) );
  nand2_1 U23711 ( .ip1(n21185), .ip2(n20959), .op(n20934) );
  nand2_1 U23712 ( .ip1(n21186), .ip2(\pipeline/csr/mcause[31] ), .op(n20932)
         );
  nand3_1 U23713 ( .ip1(n20934), .ip2(n20933), .ip3(n20932), .op(n8736) );
  nand2_1 U23714 ( .ip1(n22008), .ip2(n20959), .op(n20938) );
  xor2_1 U23715 ( .ip1(n20935), .ip2(\pipeline/csr/mtime_full [31]), .op(
        n20936) );
  nand2_1 U23716 ( .ip1(n20936), .ip2(n22009), .op(n20937) );
  nand2_1 U23717 ( .ip1(n20938), .ip2(n20937), .op(\pipeline/csr/N2112 ) );
  nand2_1 U23718 ( .ip1(n22013), .ip2(\pipeline/csr/mscratch [31]), .op(n20940) );
  nand2_1 U23719 ( .ip1(n22014), .ip2(n20959), .op(n20939) );
  nand2_1 U23720 ( .ip1(n20940), .ip2(n20939), .op(n9897) );
  nand2_1 U23721 ( .ip1(n22372), .ip2(\pipeline/csr/from_host [31]), .op(
        n20942) );
  nand2_1 U23722 ( .ip1(n22373), .ip2(n20959), .op(n20941) );
  nand2_1 U23723 ( .ip1(n20942), .ip2(n20941), .op(n9929) );
  nand2_1 U23724 ( .ip1(n22378), .ip2(n20959), .op(n20944) );
  nand2_1 U23725 ( .ip1(n22376), .ip2(\pipeline/csr/to_host [31]), .op(n20943)
         );
  nand2_1 U23726 ( .ip1(n20944), .ip2(n20943), .op(n8741) );
  inv_1 U23727 ( .ip(n20945), .op(n20946) );
  nor2_1 U23728 ( .ip1(\pipeline/csr/cycle_full [31]), .ip2(n20946), .op(
        n20948) );
  nor3_1 U23729 ( .ip1(n22289), .ip2(n20948), .ip3(n21215), .op(n20947) );
  not_ab_or_c_or_d U23730 ( .ip1(n21076), .ip2(n20959), .ip3(n21120), .ip4(
        n20947), .op(n20951) );
  nor2_1 U23731 ( .ip1(n20948), .ip2(n22289), .op(n20949) );
  nor2_1 U23732 ( .ip1(n22254), .ip2(n20949), .op(n20950) );
  nor2_1 U23733 ( .ip1(n20951), .ip2(n20950), .op(\pipeline/csr/N1904 ) );
  nand2_1 U23734 ( .ip1(n22363), .ip2(\pipeline/csr/mtimecmp [31]), .op(n20953) );
  nand2_1 U23735 ( .ip1(n22365), .ip2(n20959), .op(n20952) );
  nand2_1 U23736 ( .ip1(n20953), .ip2(n20952), .op(n9991) );
  mux2_1 U23737 ( .ip1(n20956), .ip2(\pipeline/csr/instret_full [31]), .s(
        n20954), .op(n20955) );
  nor2_1 U23738 ( .ip1(n21005), .ip2(n20955), .op(n20958) );
  nor2_1 U23739 ( .ip1(n20990), .ip2(n20956), .op(n20957) );
  ab_or_c_or_d U23740 ( .ip1(n21019), .ip2(n20959), .ip3(n20958), .ip4(n20957), 
        .op(n10107) );
  nand2_1 U23741 ( .ip1(\pipeline/csr/mie [31]), .ip2(n22356), .op(n20961) );
  nand2_1 U23742 ( .ip1(n22357), .ip2(n20959), .op(n20960) );
  nand2_1 U23743 ( .ip1(n20961), .ip2(n20960), .op(n10029) );
  nand2_1 U23744 ( .ip1(\pipeline/csr/mie [3]), .ip2(n22356), .op(n20963) );
  nand2_1 U23745 ( .ip1(n22357), .ip2(n21223), .op(n20962) );
  nand2_1 U23746 ( .ip1(n20963), .ip2(n20962), .op(n10057) );
  nor2_1 U23747 ( .ip1(\pipeline/csr/priv_stack_0 ), .ip2(n20972), .op(n20968)
         );
  nand2_1 U23748 ( .ip1(n20965), .ip2(n20964), .op(n22036) );
  and2_1 U23749 ( .ip1(n22036), .ip2(n20966), .op(n21083) );
  inv_1 U23750 ( .ip(n21083), .op(n20967) );
  nor2_1 U23751 ( .ip1(n20968), .ip2(n20967), .op(n20971) );
  nor2_1 U23752 ( .ip1(n21089), .ip2(n22036), .op(n21091) );
  inv_1 U23753 ( .ip(n21091), .op(n20969) );
  nor2_1 U23754 ( .ip1(n22268), .ip2(n20969), .op(n20970) );
  nor2_1 U23755 ( .ip1(n20971), .ip2(n20970), .op(n20974) );
  nand3_1 U23756 ( .ip1(n20972), .ip2(n21083), .ip3(n21088), .op(n22037) );
  nor2_1 U23757 ( .ip1(\pipeline/csr/priv_stack [3]), .ip2(n22037), .op(n20973) );
  nor2_1 U23758 ( .ip1(n20974), .ip2(n20973), .op(n10024) );
  nand2_1 U23759 ( .ip1(n21091), .ip2(n22377), .op(n20978) );
  nand3_1 U23760 ( .ip1(n20975), .ip2(\pipeline/csr/priv_stack [3]), .ip3(
        n21083), .op(n20977) );
  inv_1 U23761 ( .ip(n22037), .op(n21084) );
  nand2_1 U23762 ( .ip1(n21084), .ip2(\pipeline/csr/priv_stack_0 ), .op(n20976) );
  nand3_1 U23763 ( .ip1(n20978), .ip2(n20977), .ip3(n20976), .op(n10027) );
  nand2_1 U23764 ( .ip1(n21193), .ip2(n22257), .op(n20979) );
  nand2_1 U23765 ( .ip1(n20980), .ip2(n20979), .op(n20982) );
  nand2_1 U23766 ( .ip1(n22008), .ip2(n22377), .op(n20981) );
  nand2_1 U23767 ( .ip1(n20982), .ip2(n20981), .op(\pipeline/csr/N2081 ) );
  nand2_1 U23768 ( .ip1(n22013), .ip2(\pipeline/csr/mscratch [0]), .op(n20984)
         );
  nand2_1 U23769 ( .ip1(n22014), .ip2(n22377), .op(n20983) );
  nand2_1 U23770 ( .ip1(n20984), .ip2(n20983), .op(n9928) );
  inv_1 U23771 ( .ip(n21145), .op(n22022) );
  inv_1 U23772 ( .ip(\pipeline/csr/cycle_full [0]), .op(n20985) );
  nand2_1 U23773 ( .ip1(n22022), .ip2(n20985), .op(n20987) );
  nand2_1 U23774 ( .ip1(n22021), .ip2(n22377), .op(n20986) );
  nand2_1 U23775 ( .ip1(n20987), .ip2(n20986), .op(\pipeline/csr/N1873 ) );
  nand2_1 U23776 ( .ip1(n22363), .ip2(\pipeline/csr/mtimecmp [0]), .op(n20989)
         );
  nand2_1 U23777 ( .ip1(n22365), .ip2(n22377), .op(n20988) );
  nand2_1 U23778 ( .ip1(n20989), .ip2(n20988), .op(n10022) );
  mux2_1 U23779 ( .ip1(n21005), .ip2(n20990), .s(
        \pipeline/csr/instret_full [0]), .op(n20992) );
  nand2_1 U23780 ( .ip1(n21019), .ip2(n22377), .op(n20991) );
  nand2_1 U23781 ( .ip1(n20992), .ip2(n20991), .op(n10138) );
  nor2_1 U23782 ( .ip1(n22261), .ip2(n21001), .op(n20996) );
  inv_1 U23783 ( .ip(n20997), .op(n20994) );
  nor2_1 U23784 ( .ip1(\pipeline/csr/instret_full [0]), .ip2(
        \pipeline/csr/instret_full [1]), .op(n20993) );
  nor3_1 U23785 ( .ip1(n21005), .ip2(n20994), .ip3(n20993), .op(n20995) );
  ab_or_c_or_d U23786 ( .ip1(\pipeline/csr/instret_full [1]), .ip2(n21016), 
        .ip3(n20996), .ip4(n20995), .op(n10137) );
  inv_1 U23787 ( .ip(n22351), .op(n22134) );
  nor2_1 U23788 ( .ip1(n22134), .ip2(n21001), .op(n21000) );
  not_ab_or_c_or_d U23789 ( .ip1(n20998), .ip2(n20997), .ip3(n21002), .ip4(
        n21005), .op(n20999) );
  ab_or_c_or_d U23790 ( .ip1(\pipeline/csr/instret_full [2]), .ip2(n21016), 
        .ip3(n21000), .ip4(n20999), .op(n10136) );
  nor2_1 U23791 ( .ip1(n22268), .ip2(n21001), .op(n21007) );
  inv_1 U23792 ( .ip(n21008), .op(n21004) );
  nor2_1 U23793 ( .ip1(\pipeline/csr/instret_full [3]), .ip2(n21002), .op(
        n21003) );
  nor3_1 U23794 ( .ip1(n21005), .ip2(n21004), .ip3(n21003), .op(n21006) );
  ab_or_c_or_d U23795 ( .ip1(n21016), .ip2(\pipeline/csr/instret_full [3]), 
        .ip3(n21007), .ip4(n21006), .op(n10135) );
  mux2_1 U23796 ( .ip1(\pipeline/csr/instret_full [4]), .ip2(n21009), .s(
        n21008), .op(n21014) );
  inv_1 U23797 ( .ip(n21010), .op(n21011) );
  nor2_1 U23798 ( .ip1(n21012), .ip2(n21011), .op(n21013) );
  nor2_1 U23799 ( .ip1(n21014), .ip2(n21013), .op(n21015) );
  or2_1 U23800 ( .ip1(\pipeline/csr/instret_full [4]), .ip2(n21015), .op(
        n21018) );
  or2_1 U23801 ( .ip1(n21016), .ip2(n21015), .op(n21017) );
  nand2_1 U23802 ( .ip1(n21018), .ip2(n21017), .op(n21021) );
  nand2_1 U23803 ( .ip1(n21019), .ip2(n22360), .op(n21020) );
  nand2_1 U23804 ( .ip1(n21021), .ip2(n21020), .op(n10134) );
  nand2_1 U23805 ( .ip1(n22314), .ip2(n22360), .op(n21024) );
  or2_1 U23806 ( .ip1(\pipeline/csr/cycle_full [36]), .ip2(n21226), .op(n21022) );
  nand3_1 U23807 ( .ip1(n21070), .ip2(n21022), .ip3(n22316), .op(n21023) );
  nand2_1 U23808 ( .ip1(n21024), .ip2(n21023), .op(\pipeline/csr/N1909 ) );
  nand2_1 U23809 ( .ip1(n21091), .ip2(n22360), .op(n21027) );
  nand3_1 U23810 ( .ip1(\pipeline/prv [0]), .ip2(n21083), .ip3(n21082), .op(
        n21026) );
  nand2_1 U23811 ( .ip1(n21084), .ip2(\pipeline/csr/priv_stack [4]), .op(
        n21025) );
  nand3_1 U23812 ( .ip1(n21027), .ip2(n21026), .ip3(n21025), .op(n10023) );
  mux2_1 U23813 ( .ip1(\pipeline/csr_rdata_WB [4]), .ip2(n21028), .s(n19498), 
        .op(n8802) );
  mux2_1 U23814 ( .ip1(dmem_haddr[3]), .ip2(\pipeline/alu_out_WB [3]), .s(
        n21582), .op(n8729) );
  nor2_1 U23815 ( .ip1(n21223), .ip2(n21029), .op(n21034) );
  inv_1 U23816 ( .ip(\pipeline/csr/mtvec [3]), .op(n21030) );
  nor2_1 U23817 ( .ip1(n21089), .ip2(n21030), .op(n21031) );
  nor2_1 U23818 ( .ip1(n21032), .ip2(n21031), .op(n21033) );
  nor2_1 U23819 ( .ip1(n21034), .ip2(n21033), .op(n9989) );
  nor2_1 U23820 ( .ip1(n21036), .ip2(n21035), .op(n21038) );
  xor2_1 U23821 ( .ip1(n21038), .ip2(n21037), .op(imem_haddr[5]) );
  nand2_1 U23822 ( .ip1(n21995), .ip2(imem_haddr[5]), .op(n21040) );
  nand2_1 U23823 ( .ip1(\pipeline/PC_IF [5]), .ip2(n21996), .op(n21039) );
  nand2_1 U23824 ( .ip1(n21040), .ip2(n21039), .op(n8480) );
  nand2_1 U23825 ( .ip1(\pipeline/PC_IF [5]), .ip2(n21988), .op(n21042) );
  nand2_1 U23826 ( .ip1(\pipeline/PC_DX [5]), .ip2(n21999), .op(n21041) );
  nand2_1 U23827 ( .ip1(n21042), .ip2(n21041), .op(n8479) );
  mux2_1 U23828 ( .ip1(\pipeline/PC_WB [5]), .ip2(\pipeline/PC_DX [5]), .s(
        n17429), .op(n8898) );
  nand2_1 U23829 ( .ip1(n21043), .ip2(n22145), .op(n21049) );
  xor2_1 U23830 ( .ip1(\pipeline/PC_WB [5]), .ip2(n21044), .op(n21045) );
  nand2_1 U23831 ( .ip1(n21046), .ip2(n21045), .op(n21048) );
  nand2_1 U23832 ( .ip1(\pipeline/epc [5]), .ip2(n21174), .op(n21047) );
  nand3_1 U23833 ( .ip1(n21049), .ip2(n21048), .ip3(n21047), .op(n8866) );
  inv_1 U23834 ( .ip(n22145), .op(n21067) );
  nor2_1 U23835 ( .ip1(n21067), .ip2(n22267), .op(n21054) );
  not_ab_or_c_or_d U23836 ( .ip1(n21052), .ip2(n21051), .ip3(n21050), .ip4(
        n22276), .op(n21053) );
  or2_1 U23837 ( .ip1(n21054), .ip2(n21053), .op(\pipeline/csr/N1974 ) );
  inv_1 U23838 ( .ip(n21055), .op(n21056) );
  nor2_1 U23839 ( .ip1(\pipeline/csr/time_full [5]), .ip2(n21056), .op(n21059)
         );
  nor3_1 U23840 ( .ip1(n21177), .ip2(n21058), .ip3(n21059), .op(n21057) );
  not_ab_or_c_or_d U23841 ( .ip1(n21179), .ip2(n22145), .ip3(n21120), .ip4(
        n21057), .op(n21062) );
  nor2_1 U23842 ( .ip1(n21059), .ip2(n21058), .op(n21060) );
  nor2_1 U23843 ( .ip1(n21198), .ip2(n21060), .op(n21061) );
  nor2_1 U23844 ( .ip1(n21062), .ip2(n21061), .op(\pipeline/csr/N1942 ) );
  nand2_1 U23845 ( .ip1(n22008), .ip2(n22145), .op(n21066) );
  xor2_1 U23846 ( .ip1(\pipeline/csr/mtime_full [5]), .ip2(n21063), .op(n21064) );
  nand2_1 U23847 ( .ip1(n21064), .ip2(n22009), .op(n21065) );
  nand2_1 U23848 ( .ip1(n21066), .ip2(n21065), .op(\pipeline/csr/N2086 ) );
  nor2_1 U23849 ( .ip1(n21067), .ip2(n22305), .op(n21072) );
  not_ab_or_c_or_d U23850 ( .ip1(n21070), .ip2(n21069), .ip3(n21068), .ip4(
        n22308), .op(n21071) );
  or2_1 U23851 ( .ip1(n21072), .ip2(n21071), .op(\pipeline/csr/N1910 ) );
  inv_1 U23852 ( .ip(n21073), .op(n21074) );
  nor2_1 U23853 ( .ip1(\pipeline/csr/cycle_full [5]), .ip2(n21074), .op(n21078) );
  nor3_1 U23854 ( .ip1(n21077), .ip2(n21078), .ip3(n21215), .op(n21075) );
  not_ab_or_c_or_d U23855 ( .ip1(n21076), .ip2(n22145), .ip3(n21217), .ip4(
        n21075), .op(n21081) );
  nor2_1 U23856 ( .ip1(n21078), .ip2(n21077), .op(n21079) );
  nor2_1 U23857 ( .ip1(n22254), .ip2(n21079), .op(n21080) );
  nor2_1 U23858 ( .ip1(n21081), .ip2(n21080), .op(\pipeline/csr/N1878 ) );
  nand2_1 U23859 ( .ip1(n21091), .ip2(n22145), .op(n21087) );
  nand3_1 U23860 ( .ip1(\pipeline/prv [1]), .ip2(n21083), .ip3(n21082), .op(
        n21086) );
  nand2_1 U23861 ( .ip1(n21084), .ip2(\pipeline/csr/priv_stack [5]), .op(
        n21085) );
  nand3_1 U23862 ( .ip1(n21087), .ip2(n21086), .ip3(n21085), .op(n10028) );
  nor2_1 U23863 ( .ip1(n21089), .ip2(n21088), .op(n21090) );
  nor2_1 U23864 ( .ip1(n21091), .ip2(n21090), .op(n22034) );
  nor2_1 U23865 ( .ip1(n22134), .ip2(n22036), .op(n21092) );
  not_ab_or_c_or_d U23866 ( .ip1(\pipeline/csr/priv_stack [5]), .ip2(n22036), 
        .ip3(n22034), .ip4(n21092), .op(n21094) );
  nor2_1 U23867 ( .ip1(\pipeline/prv [1]), .ip2(n22037), .op(n21093) );
  nor2_1 U23868 ( .ip1(n21094), .ip2(n21093), .op(n10025) );
  nand2_1 U23869 ( .ip1(\pipeline/ctrl/prev_ex_code_WB [1]), .ip2(n19505), 
        .op(n21101) );
  nand2_1 U23870 ( .ip1(\pipeline/prv [1]), .ip2(n21095), .op(n21096) );
  nand2_1 U23871 ( .ip1(n21097), .ip2(n21096), .op(n21098) );
  nand2_1 U23872 ( .ip1(n21099), .ip2(n21098), .op(n21100) );
  nand2_1 U23873 ( .ip1(n21101), .ip2(n21100), .op(n8737) );
  mux2_1 U23874 ( .ip1(dmem_haddr[2]), .ip2(\pipeline/alu_out_WB [2]), .s(
        n19505), .op(n8730) );
  nand2_1 U23875 ( .ip1(n22282), .ip2(n22351), .op(n21104) );
  or2_1 U23876 ( .ip1(\pipeline/csr/time_full [34]), .ip2(n22262), .op(n21102)
         );
  nand3_1 U23877 ( .ip1(n21102), .ip2(n22270), .ip3(n22284), .op(n21103) );
  nand2_1 U23878 ( .ip1(n21104), .ip2(n21103), .op(\pipeline/csr/N1971 ) );
  nor2_1 U23879 ( .ip1(n22261), .ip2(n21110), .op(n21109) );
  inv_1 U23880 ( .ip(n21113), .op(n21107) );
  nor2_1 U23881 ( .ip1(\pipeline/csr/instret_full [33]), .ip2(n21105), .op(
        n21106) );
  nor3_1 U23882 ( .ip1(n21111), .ip2(n21107), .ip3(n21106), .op(n21108) );
  ab_or_c_or_d U23883 ( .ip1(\pipeline/csr/instret_full [33]), .ip2(n21117), 
        .ip3(n21109), .ip4(n21108), .op(n10105) );
  nor2_1 U23884 ( .ip1(n22134), .ip2(n21110), .op(n21116) );
  not_ab_or_c_or_d U23885 ( .ip1(n21114), .ip2(n21113), .ip3(n21112), .ip4(
        n21111), .op(n21115) );
  ab_or_c_or_d U23886 ( .ip1(\pipeline/csr/instret_full [34]), .ip2(n21117), 
        .ip3(n21116), .ip4(n21115), .op(n10104) );
  nand2_1 U23887 ( .ip1(\pipeline/csr/time_full [1]), .ip2(
        \pipeline/csr/time_full [0]), .op(n21118) );
  xor2_1 U23888 ( .ip1(\pipeline/csr/time_full [2]), .ip2(n21118), .op(n21121)
         );
  nor2_1 U23889 ( .ip1(n21177), .ip2(n21121), .op(n21119) );
  not_ab_or_c_or_d U23890 ( .ip1(n21179), .ip2(n22351), .ip3(n21120), .ip4(
        n21119), .op(n21124) );
  inv_1 U23891 ( .ip(n21121), .op(n21122) );
  nor2_1 U23892 ( .ip1(n21198), .ip2(n21122), .op(n21123) );
  nor2_1 U23893 ( .ip1(n21124), .ip2(n21123), .op(\pipeline/csr/N1939 ) );
  nand2_1 U23894 ( .ip1(n22351), .ip2(n21185), .op(n21130) );
  inv_1 U23895 ( .ip(\pipeline/csr/mecode [2]), .op(n21126) );
  nor2_1 U23896 ( .ip1(n21126), .ip2(n21125), .op(n21127) );
  nor2_1 U23897 ( .ip1(n21128), .ip2(n21127), .op(n21129) );
  nand2_1 U23898 ( .ip1(n21130), .ip2(n21129), .op(n8733) );
  nor2_1 U23899 ( .ip1(n22134), .ip2(n21131), .op(n21136) );
  nand2_1 U23900 ( .ip1(\pipeline/csr/mtime_full [1]), .ip2(
        \pipeline/csr/mtime_full [0]), .op(n21132) );
  xor2_1 U23901 ( .ip1(\pipeline/csr/mtime_full [2]), .ip2(n21132), .op(n21133) );
  nor2_1 U23902 ( .ip1(n21134), .ip2(n21133), .op(n21135) );
  or2_1 U23903 ( .ip1(n21136), .ip2(n21135), .op(\pipeline/csr/N2083 ) );
  nand2_1 U23904 ( .ip1(\pipeline/csr/mscratch [2]), .ip2(n22013), .op(n21138)
         );
  nand2_1 U23905 ( .ip1(n22014), .ip2(n22351), .op(n21137) );
  nand2_1 U23906 ( .ip1(n21138), .ip2(n21137), .op(n9926) );
  nand2_1 U23907 ( .ip1(\pipeline/csr/from_host [2]), .ip2(n22372), .op(n21140) );
  nand2_1 U23908 ( .ip1(n22373), .ip2(n22351), .op(n21139) );
  nand2_1 U23909 ( .ip1(n21140), .ip2(n21139), .op(n9958) );
  nand2_1 U23910 ( .ip1(n22378), .ip2(n22351), .op(n21142) );
  nand2_1 U23911 ( .ip1(\pipeline/csr/to_host [2]), .ip2(n22376), .op(n21141)
         );
  nand2_1 U23912 ( .ip1(n21142), .ip2(n21141), .op(n8770) );
  nand2_1 U23913 ( .ip1(n22021), .ip2(n22351), .op(n21147) );
  nand2_1 U23914 ( .ip1(\pipeline/csr/cycle_full [1]), .ip2(
        \pipeline/csr/cycle_full [0]), .op(n21143) );
  xor2_1 U23915 ( .ip1(\pipeline/csr/cycle_full [2]), .ip2(n21143), .op(n21144) );
  or2_1 U23916 ( .ip1(n21145), .ip2(n21144), .op(n21146) );
  nand2_1 U23917 ( .ip1(n21147), .ip2(n21146), .op(\pipeline/csr/N1875 ) );
  nand2_1 U23918 ( .ip1(\pipeline/csr/mtimecmp [2]), .ip2(n22363), .op(n21149)
         );
  nand2_1 U23919 ( .ip1(n22365), .ip2(n22351), .op(n21148) );
  nand2_1 U23920 ( .ip1(n21149), .ip2(n21148), .op(n10020) );
  mux2_1 U23921 ( .ip1(\pipeline/csr_rdata_WB [2]), .ip2(n21150), .s(n19498), 
        .op(n8804) );
  inv_1 U23922 ( .ip(dmem_rdata[26]), .op(n21151) );
  nor2_1 U23923 ( .ip1(n21233), .ip2(n21151), .op(n21154) );
  inv_1 U23924 ( .ip(dmem_rdata[10]), .op(n21152) );
  nor2_1 U23925 ( .ip1(n21235), .ip2(n21152), .op(n21153) );
  not_ab_or_c_or_d U23926 ( .ip1(n21238), .ip2(dmem_rdata[2]), .ip3(n21154), 
        .ip4(n21153), .op(n21158) );
  nand2_1 U23927 ( .ip1(n21155), .ip2(n21583), .op(n21157) );
  nand2_1 U23928 ( .ip1(n21240), .ip2(dmem_rdata[18]), .op(n21156) );
  nand3_1 U23929 ( .ip1(n21158), .ip2(n21157), .ip3(n21156), .op(n21159) );
  mux2_1 U23930 ( .ip1(\pipeline/regfile/data[22][2] ), .ip2(n21159), .s(
        n21589), .op(n9222) );
  mux2_1 U23931 ( .ip1(\pipeline/regfile/data[28][2] ), .ip2(n21159), .s(
        n21590), .op(n9030) );
  mux2_1 U23932 ( .ip1(\pipeline/regfile/data[12][2] ), .ip2(n21159), .s(
        n21591), .op(n9542) );
  mux2_1 U23933 ( .ip1(\pipeline/regfile/data[19][2] ), .ip2(n21159), .s(
        n21592), .op(n9318) );
  mux2_1 U23934 ( .ip1(\pipeline/regfile/data[11][2] ), .ip2(n21159), .s(
        n21593), .op(n9574) );
  mux2_1 U23935 ( .ip1(\pipeline/regfile/data[30][2] ), .ip2(n21159), .s(
        n21594), .op(n8966) );
  mux2_1 U23936 ( .ip1(\pipeline/regfile/data[18][2] ), .ip2(n21159), .s(
        n21595), .op(n9350) );
  mux2_1 U23937 ( .ip1(\pipeline/regfile/data[23][2] ), .ip2(n21159), .s(
        n21596), .op(n9190) );
  mux2_1 U23938 ( .ip1(\pipeline/regfile/data[6][2] ), .ip2(n21159), .s(n21597), .op(n9734) );
  mux2_1 U23939 ( .ip1(\pipeline/regfile/data[5][2] ), .ip2(n21159), .s(n21598), .op(n9766) );
  mux2_1 U23940 ( .ip1(\pipeline/regfile/data[3][2] ), .ip2(n21159), .s(n21599), .op(n9830) );
  mux2_1 U23941 ( .ip1(\pipeline/regfile/data[13][2] ), .ip2(n21159), .s(
        n21600), .op(n9510) );
  mux2_1 U23942 ( .ip1(\pipeline/regfile/data[20][2] ), .ip2(n21159), .s(
        n21601), .op(n9286) );
  mux2_1 U23943 ( .ip1(\pipeline/regfile/data[25][2] ), .ip2(n21159), .s(
        n21602), .op(n9126) );
  mux2_1 U23944 ( .ip1(\pipeline/regfile/data[24][2] ), .ip2(n21159), .s(
        n21603), .op(n9158) );
  mux2_1 U23945 ( .ip1(\pipeline/regfile/data[14][2] ), .ip2(n21159), .s(
        n21604), .op(n9478) );
  mux2_1 U23946 ( .ip1(\pipeline/regfile/data[4][2] ), .ip2(n21159), .s(n21605), .op(n9798) );
  mux2_1 U23947 ( .ip1(\pipeline/regfile/data[31][2] ), .ip2(n21159), .s(
        n21606), .op(n8934) );
  mux2_1 U23948 ( .ip1(\pipeline/regfile/data[26][2] ), .ip2(n21159), .s(
        n21607), .op(n9094) );
  mux2_1 U23949 ( .ip1(\pipeline/regfile/data[16][2] ), .ip2(n21159), .s(
        n21608), .op(n9414) );
  mux2_1 U23950 ( .ip1(\pipeline/regfile/data[9][2] ), .ip2(n21159), .s(n21609), .op(n9638) );
  mux2_1 U23951 ( .ip1(\pipeline/regfile/data[2][2] ), .ip2(n21159), .s(n21610), .op(n9862) );
  mux2_1 U23952 ( .ip1(\pipeline/regfile/data[1][2] ), .ip2(n21159), .s(n21611), .op(n9894) );
  mux2_1 U23953 ( .ip1(\pipeline/regfile/data[27][2] ), .ip2(n21159), .s(
        n21612), .op(n9062) );
  mux2_1 U23954 ( .ip1(\pipeline/regfile/data[15][2] ), .ip2(n21159), .s(
        n21613), .op(n9446) );
  mux2_1 U23955 ( .ip1(\pipeline/regfile/data[7][2] ), .ip2(n21159), .s(n21614), .op(n9702) );
  mux2_1 U23956 ( .ip1(\pipeline/regfile/data[21][2] ), .ip2(n21159), .s(
        n21615), .op(n9254) );
  mux2_1 U23957 ( .ip1(\pipeline/regfile/data[17][2] ), .ip2(n21159), .s(
        n21616), .op(n9382) );
  mux2_1 U23958 ( .ip1(\pipeline/regfile/data[8][2] ), .ip2(n21159), .s(n21617), .op(n9670) );
  mux2_1 U23959 ( .ip1(\pipeline/regfile/data[10][2] ), .ip2(n21159), .s(
        n21618), .op(n9606) );
  mux2_1 U23960 ( .ip1(\pipeline/regfile/data[29][2] ), .ip2(n21159), .s(
        n21619), .op(n8998) );
  nor2_1 U23961 ( .ip1(n21161), .ip2(n21160), .op(n21163) );
  xor2_1 U23962 ( .ip1(n21163), .ip2(n21162), .op(imem_haddr[3]) );
  nand2_1 U23963 ( .ip1(n21995), .ip2(imem_haddr[3]), .op(n21165) );
  nand2_1 U23964 ( .ip1(\pipeline/PC_IF [3]), .ip2(n21996), .op(n21164) );
  nand2_1 U23965 ( .ip1(n21165), .ip2(n21164), .op(n8484) );
  nand2_1 U23966 ( .ip1(\pipeline/PC_IF [3]), .ip2(n22048), .op(n21167) );
  nand2_1 U23967 ( .ip1(\pipeline/PC_DX [3]), .ip2(n21999), .op(n21166) );
  nand2_1 U23968 ( .ip1(n21167), .ip2(n21166), .op(n8483) );
  mux2_1 U23969 ( .ip1(\pipeline/PC_WB [3]), .ip2(\pipeline/PC_DX [3]), .s(
        n17777), .op(n8900) );
  nor2_1 U23970 ( .ip1(n22268), .ip2(n21168), .op(n21173) );
  xor2_1 U23971 ( .ip1(\pipeline/PC_WB [3]), .ip2(n21169), .op(n21170) );
  nor2_1 U23972 ( .ip1(n21171), .ip2(n21170), .op(n21172) );
  ab_or_c_or_d U23973 ( .ip1(n21174), .ip2(\pipeline/epc [3]), .ip3(n21173), 
        .ip4(n21172), .op(n8868) );
  inv_1 U23974 ( .ip(n21175), .op(n21176) );
  nor2_1 U23975 ( .ip1(\pipeline/csr/time_full [3]), .ip2(n21176), .op(n21181)
         );
  nor3_1 U23976 ( .ip1(n21177), .ip2(n21180), .ip3(n21181), .op(n21178) );
  not_ab_or_c_or_d U23977 ( .ip1(n21179), .ip2(n21223), .ip3(n21217), .ip4(
        n21178), .op(n21184) );
  nor2_1 U23978 ( .ip1(n21181), .ip2(n21180), .op(n21182) );
  nor2_1 U23979 ( .ip1(n22254), .ip2(n21182), .op(n21183) );
  nor2_1 U23980 ( .ip1(n21184), .ip2(n21183), .op(\pipeline/csr/N1940 ) );
  nand2_1 U23981 ( .ip1(n21185), .ip2(n21223), .op(n21190) );
  nand2_1 U23982 ( .ip1(\pipeline/csr/mecode [3]), .ip2(n21186), .op(n21189)
         );
  nand2_1 U23983 ( .ip1(n21187), .ip2(\pipeline/ctrl/prev_ex_code_WB [3]), 
        .op(n21188) );
  nand3_1 U23984 ( .ip1(n21190), .ip2(n21189), .ip3(n21188), .op(n8732) );
  xor2_1 U23985 ( .ip1(n21192), .ip2(n21191), .op(n21196) );
  nor2_1 U23986 ( .ip1(n21193), .ip2(n21196), .op(n21194) );
  not_ab_or_c_or_d U23987 ( .ip1(n21195), .ip2(n21223), .ip3(n21217), .ip4(
        n21194), .op(n21200) );
  inv_1 U23988 ( .ip(n21196), .op(n21197) );
  nor2_1 U23989 ( .ip1(n21198), .ip2(n21197), .op(n21199) );
  nor2_1 U23990 ( .ip1(n21200), .ip2(n21199), .op(\pipeline/csr/N2084 ) );
  nand2_1 U23991 ( .ip1(\pipeline/csr/mscratch [3]), .ip2(n22013), .op(n21202)
         );
  nand2_1 U23992 ( .ip1(n22014), .ip2(n21223), .op(n21201) );
  nand2_1 U23993 ( .ip1(n21202), .ip2(n21201), .op(n9925) );
  nand2_1 U23994 ( .ip1(\pipeline/csr/from_host [3]), .ip2(n22372), .op(n21204) );
  nand2_1 U23995 ( .ip1(n22373), .ip2(n21223), .op(n21203) );
  nand2_1 U23996 ( .ip1(n21204), .ip2(n21203), .op(n9957) );
  nand2_1 U23997 ( .ip1(n22378), .ip2(n21223), .op(n21206) );
  nand2_1 U23998 ( .ip1(\pipeline/csr/to_host [3]), .ip2(n22376), .op(n21205)
         );
  nand2_1 U23999 ( .ip1(n21206), .ip2(n21205), .op(n8769) );
  xor2_1 U24000 ( .ip1(\pipeline/csr/mtime_full [35]), .ip2(n22135), .op(
        n21207) );
  nand2_1 U24001 ( .ip1(n18449), .ip2(n21207), .op(n21212) );
  nand2_1 U24002 ( .ip1(n21208), .ip2(n21223), .op(n21209) );
  or2_1 U24003 ( .ip1(n21210), .ip2(n21209), .op(n21211) );
  nand2_1 U24004 ( .ip1(n21212), .ip2(n21211), .op(\pipeline/csr/N2116 ) );
  inv_1 U24005 ( .ip(n21213), .op(n21214) );
  nor2_1 U24006 ( .ip1(\pipeline/csr/cycle_full [3]), .ip2(n21214), .op(n21219) );
  nor3_1 U24007 ( .ip1(n21218), .ip2(n21219), .ip3(n21215), .op(n21216) );
  not_ab_or_c_or_d U24008 ( .ip1(n21076), .ip2(n21223), .ip3(n21217), .ip4(
        n21216), .op(n21222) );
  nor2_1 U24009 ( .ip1(n21219), .ip2(n21218), .op(n21220) );
  nor2_1 U24010 ( .ip1(n22254), .ip2(n21220), .op(n21221) );
  nor2_1 U24011 ( .ip1(n21222), .ip2(n21221), .op(\pipeline/csr/N1876 ) );
  nand2_1 U24012 ( .ip1(\pipeline/csr/mtimecmp [3]), .ip2(n22363), .op(n21225)
         );
  nand2_1 U24013 ( .ip1(n22365), .ip2(n21223), .op(n21224) );
  nand2_1 U24014 ( .ip1(n21225), .ip2(n21224), .op(n10019) );
  nor2_1 U24015 ( .ip1(n22268), .ip2(n22305), .op(n21229) );
  not_ab_or_c_or_d U24016 ( .ip1(n22296), .ip2(n21227), .ip3(n21226), .ip4(
        n22308), .op(n21228) );
  or2_1 U24017 ( .ip1(n21229), .ip2(n21228), .op(\pipeline/csr/N1908 ) );
  nor2_1 U24018 ( .ip1(\pipeline/csr/mip_3 ), .ip2(n21231), .op(n21230) );
  not_ab_or_c_or_d U24019 ( .ip1(n22268), .ip2(n21231), .ip3(htif_reset), 
        .ip4(n21230), .op(n10074) );
  mux2_1 U24020 ( .ip1(dmem_haddr[1]), .ip2(\pipeline/alu_out_WB [1]), .s(
        n21582), .op(n8731) );
  inv_1 U24021 ( .ip(dmem_rdata[24]), .op(n21232) );
  nor2_1 U24022 ( .ip1(n21233), .ip2(n21232), .op(n21237) );
  inv_1 U24023 ( .ip(dmem_rdata[8]), .op(n21234) );
  nor2_1 U24024 ( .ip1(n21235), .ip2(n21234), .op(n21236) );
  not_ab_or_c_or_d U24025 ( .ip1(n21238), .ip2(dmem_rdata[0]), .ip3(n21237), 
        .ip4(n21236), .op(n21243) );
  nand2_1 U24026 ( .ip1(n21239), .ip2(n21583), .op(n21242) );
  nand2_1 U24027 ( .ip1(n21240), .ip2(dmem_rdata[16]), .op(n21241) );
  nand3_1 U24028 ( .ip1(n21243), .ip2(n21242), .ip3(n21241), .op(n21244) );
  mux2_1 U24029 ( .ip1(\pipeline/regfile/data[22][0] ), .ip2(n21244), .s(
        n21589), .op(n9224) );
  mux2_1 U24030 ( .ip1(\pipeline/regfile/data[28][0] ), .ip2(n21244), .s(
        n21590), .op(n9032) );
  mux2_1 U24031 ( .ip1(\pipeline/regfile/data[12][0] ), .ip2(n21244), .s(
        n21591), .op(n9544) );
  mux2_1 U24032 ( .ip1(\pipeline/regfile/data[19][0] ), .ip2(n21244), .s(
        n21592), .op(n9320) );
  mux2_1 U24033 ( .ip1(\pipeline/regfile/data[11][0] ), .ip2(n21244), .s(
        n21593), .op(n9576) );
  mux2_1 U24034 ( .ip1(\pipeline/regfile/data[30][0] ), .ip2(n21244), .s(
        n21594), .op(n8968) );
  mux2_1 U24035 ( .ip1(\pipeline/regfile/data[18][0] ), .ip2(n21244), .s(
        n21595), .op(n9352) );
  mux2_1 U24036 ( .ip1(\pipeline/regfile/data[23][0] ), .ip2(n21244), .s(
        n21596), .op(n9192) );
  mux2_1 U24037 ( .ip1(\pipeline/regfile/data[6][0] ), .ip2(n21244), .s(n21597), .op(n9736) );
  mux2_1 U24038 ( .ip1(\pipeline/regfile/data[5][0] ), .ip2(n21244), .s(n21598), .op(n9768) );
  mux2_1 U24039 ( .ip1(\pipeline/regfile/data[3][0] ), .ip2(n21244), .s(n21599), .op(n9832) );
  mux2_1 U24040 ( .ip1(\pipeline/regfile/data[13][0] ), .ip2(n21244), .s(
        n21600), .op(n9512) );
  mux2_1 U24041 ( .ip1(\pipeline/regfile/data[20][0] ), .ip2(n21244), .s(
        n21601), .op(n9288) );
  mux2_1 U24042 ( .ip1(\pipeline/regfile/data[25][0] ), .ip2(n21244), .s(
        n21602), .op(n9128) );
  mux2_1 U24043 ( .ip1(\pipeline/regfile/data[24][0] ), .ip2(n21244), .s(
        n21603), .op(n9160) );
  mux2_1 U24044 ( .ip1(\pipeline/regfile/data[14][0] ), .ip2(n21244), .s(
        n21604), .op(n9480) );
  mux2_1 U24045 ( .ip1(\pipeline/regfile/data[4][0] ), .ip2(n21244), .s(n21605), .op(n9800) );
  mux2_1 U24046 ( .ip1(\pipeline/regfile/data[31][0] ), .ip2(n21244), .s(
        n21606), .op(n8936) );
  mux2_1 U24047 ( .ip1(\pipeline/regfile/data[26][0] ), .ip2(n21244), .s(
        n21607), .op(n9096) );
  mux2_1 U24048 ( .ip1(\pipeline/regfile/data[16][0] ), .ip2(n21244), .s(
        n21608), .op(n9416) );
  mux2_1 U24049 ( .ip1(\pipeline/regfile/data[9][0] ), .ip2(n21244), .s(n21609), .op(n9640) );
  mux2_1 U24050 ( .ip1(\pipeline/regfile/data[2][0] ), .ip2(n21244), .s(n21610), .op(n9864) );
  mux2_1 U24051 ( .ip1(\pipeline/regfile/data[1][0] ), .ip2(n21244), .s(n21611), .op(n9896) );
  mux2_1 U24052 ( .ip1(\pipeline/regfile/data[27][0] ), .ip2(n21244), .s(
        n21612), .op(n9064) );
  mux2_1 U24053 ( .ip1(\pipeline/regfile/data[15][0] ), .ip2(n21244), .s(
        n21613), .op(n9448) );
  mux2_1 U24054 ( .ip1(\pipeline/regfile/data[7][0] ), .ip2(n21244), .s(n21614), .op(n9704) );
  mux2_1 U24055 ( .ip1(\pipeline/regfile/data[21][0] ), .ip2(n21244), .s(
        n21615), .op(n9256) );
  mux2_1 U24056 ( .ip1(\pipeline/regfile/data[17][0] ), .ip2(n21244), .s(
        n21616), .op(n9384) );
  mux2_1 U24057 ( .ip1(\pipeline/regfile/data[8][0] ), .ip2(n21244), .s(n21617), .op(n9672) );
  mux2_1 U24058 ( .ip1(\pipeline/regfile/data[10][0] ), .ip2(n21244), .s(
        n21618), .op(n9608) );
  mux2_1 U24059 ( .ip1(\pipeline/regfile/data[29][0] ), .ip2(n21244), .s(
        n21619), .op(n9000) );
  inv_1 U24060 ( .ip(n21245), .op(n21246) );
  nand3_1 U24061 ( .ip1(n21248), .ip2(n21247), .ip3(n21246), .op(n21252) );
  nand2_1 U24062 ( .ip1(n21440), .ip2(n21252), .op(n21249) );
  nand2_1 U24063 ( .ip1(n21250), .ip2(n21249), .op(n21270) );
  inv_1 U24064 ( .ip(n21251), .op(n21253) );
  nor3_1 U24065 ( .ip1(\pipeline/md_resp_result [1]), .ip2(n21253), .ip3(
        n21252), .op(n21269) );
  nand2_1 U24066 ( .ip1(\pipeline/md/negate_output ), .ip2(n21520), .op(n21254) );
  nor2_1 U24067 ( .ip1(n21256), .ip2(n21254), .op(n21260) );
  nor2_1 U24068 ( .ip1(n21255), .ip2(n21957), .op(n21258) );
  nor2_1 U24069 ( .ip1(n21960), .ip2(n21256), .op(n21257) );
  nor2_1 U24070 ( .ip1(n21258), .ip2(n21257), .op(n21259) );
  nor2_1 U24071 ( .ip1(n21260), .ip2(n21259), .op(n21267) );
  inv_1 U24072 ( .ip(n21263), .op(n21261) );
  nor3_1 U24073 ( .ip1(\pipeline/md/result [33]), .ip2(n21966), .ip3(n21261), 
        .op(n21265) );
  inv_1 U24074 ( .ip(\pipeline/md/result [33]), .op(n21262) );
  not_ab_or_c_or_d U24075 ( .ip1(\pipeline/md/negate_output ), .ip2(n21263), 
        .ip3(n21262), .ip4(n21967), .op(n21264) );
  nor3_1 U24076 ( .ip1(n21972), .ip2(n21265), .ip3(n21264), .op(n21266) );
  nor2_1 U24077 ( .ip1(n21267), .ip2(n21266), .op(n21268) );
  not_ab_or_c_or_d U24078 ( .ip1(\pipeline/md_resp_result [1]), .ip2(n21270), 
        .ip3(n21269), .ip4(n21268), .op(n21274) );
  nand2_1 U24079 ( .ip1(n21272), .ip2(n21271), .op(n21273) );
  nand2_1 U24080 ( .ip1(n21274), .ip2(n21273), .op(n8633) );
  mux2_1 U24081 ( .ip1(\pipeline/csr_rdata_WB [1]), .ip2(n21275), .s(n17777), 
        .op(n8805) );
  nand2_1 U24082 ( .ip1(n21427), .ip2(n21276), .op(n21285) );
  nand2_1 U24083 ( .ip1(n21280), .ip2(n21279), .op(n21324) );
  nor2_1 U24084 ( .ip1(n21278), .ip2(n21324), .op(n21318) );
  nor2_1 U24085 ( .ip1(n21281), .ip2(n21282), .op(n21283) );
  nand2_1 U24086 ( .ip1(n21318), .ip2(n21283), .op(n21302) );
  nor2_1 U24087 ( .ip1(n21277), .ip2(n21302), .op(n21284) );
  or2_1 U24088 ( .ip1(n21284), .ip2(n21414), .op(n21298) );
  nand2_1 U24089 ( .ip1(n21285), .ip2(n21298), .op(n21293) );
  not_ab_or_c_or_d U24090 ( .ip1(n21427), .ip2(n22063), .ip3(n22066), .ip4(
        n21293), .op(n21682) );
  inv_1 U24091 ( .ip(n22066), .op(n21287) );
  nor2_1 U24092 ( .ip1(n22063), .ip2(n21293), .op(n21286) );
  nor2_1 U24093 ( .ip1(n21287), .ip2(n21286), .op(n21288) );
  nor2_1 U24094 ( .ip1(n21288), .ip2(n21683), .op(n21289) );
  nor2_1 U24095 ( .ip1(n21400), .ip2(n21289), .op(n21290) );
  nor2_1 U24096 ( .ip1(n21682), .ip2(n21290), .op(n21292) );
  nor2_1 U24097 ( .ip1(n22744), .ip2(n21680), .op(n21291) );
  ab_or_c_or_d U24098 ( .ip1(n14765), .ip2(\pipeline/md/b [62]), .ip3(n21292), 
        .ip4(n21291), .op(n8422) );
  xor2_1 U24099 ( .ip1(n22063), .ip2(n21293), .op(n21294) );
  nand2_1 U24100 ( .ip1(n22042), .ip2(n21294), .op(n21297) );
  nand2_1 U24101 ( .ip1(\pipeline/md/b [61]), .ip2(n20310), .op(n21296) );
  nand2_1 U24102 ( .ip1(\pipeline/md/b [60]), .ip2(n21496), .op(n21295) );
  nand3_1 U24103 ( .ip1(n21297), .ip2(n21296), .ip3(n21295), .op(n8418) );
  nor2_1 U24104 ( .ip1(n22734), .ip2(n22665), .op(n21301) );
  xor2_1 U24105 ( .ip1(n21276), .ip2(n21298), .op(n21299) );
  nor2_1 U24106 ( .ip1(n21299), .ip2(n21683), .op(n21300) );
  ab_or_c_or_d U24107 ( .ip1(n21493), .ip2(\pipeline/md/b [59]), .ip3(n21301), 
        .ip4(n21300), .op(n8417) );
  nand2_1 U24108 ( .ip1(n21302), .ip2(n21360), .op(n21314) );
  nor2_1 U24109 ( .ip1(n21683), .ip2(n21302), .op(n21303) );
  nor2_1 U24110 ( .ip1(n21400), .ip2(n21303), .op(n21304) );
  mux2_1 U24111 ( .ip1(n21314), .ip2(n21304), .s(n21277), .op(n21307) );
  nand2_1 U24112 ( .ip1(n21493), .ip2(\pipeline/md/b [58]), .op(n21306) );
  nand2_1 U24113 ( .ip1(n21440), .ip2(\pipeline/md/b [59]), .op(n21305) );
  nand3_1 U24114 ( .ip1(n21307), .ip2(n21306), .ip3(n21305), .op(n8416) );
  nor2_1 U24115 ( .ip1(n22665), .ip2(n21308), .op(n21310) );
  nor2_1 U24116 ( .ip1(n21320), .ip2(n21680), .op(n21309) );
  nor2_1 U24117 ( .ip1(n21310), .ip2(n21309), .op(n21317) );
  nor2_1 U24118 ( .ip1(n21683), .ip2(n21324), .op(n21325) );
  nor2_1 U24119 ( .ip1(n21282), .ip2(n21278), .op(n21311) );
  nand2_1 U24120 ( .ip1(n21325), .ip2(n21311), .op(n21312) );
  and2_1 U24121 ( .ip1(n21312), .ip2(n21409), .op(n21315) );
  inv_1 U24122 ( .ip(n21281), .op(n21313) );
  mux2_1 U24123 ( .ip1(n21315), .ip2(n21314), .s(n21313), .op(n21316) );
  nand2_1 U24124 ( .ip1(n21317), .ip2(n21316), .op(n8413) );
  nor2_1 U24125 ( .ip1(n21318), .ip2(n21414), .op(n21319) );
  xor2_1 U24126 ( .ip1(n21319), .ip2(n21282), .op(n21323) );
  nor2_1 U24127 ( .ip1(n21320), .ip2(n22665), .op(n21322) );
  nor2_1 U24128 ( .ip1(n21905), .ip2(n21680), .op(n21321) );
  ab_or_c_or_d U24129 ( .ip1(n22042), .ip2(n21323), .ip3(n21322), .ip4(n21321), 
        .op(n8403) );
  nand2_1 U24130 ( .ip1(n21360), .ip2(n21324), .op(n21327) );
  nor2_1 U24131 ( .ip1(n21400), .ip2(n21325), .op(n21326) );
  mux2_1 U24132 ( .ip1(n21327), .ip2(n21326), .s(n21278), .op(n21330) );
  nand2_1 U24133 ( .ip1(\pipeline/md/b [55]), .ip2(n21496), .op(n21329) );
  nand2_1 U24134 ( .ip1(\pipeline/md/b [56]), .ip2(n20310), .op(n21328) );
  nand3_1 U24135 ( .ip1(n21330), .ip2(n21329), .ip3(n21328), .op(n8402) );
  nand2_1 U24136 ( .ip1(n21427), .ip2(n21331), .op(n21332) );
  xor2_1 U24137 ( .ip1(n22086), .ip2(n21332), .op(n21333) );
  nor2_1 U24138 ( .ip1(n21333), .ip2(n21683), .op(n21335) );
  nor2_1 U24139 ( .ip1(n22680), .ip2(n21680), .op(n21334) );
  ab_or_c_or_d U24140 ( .ip1(n14765), .ip2(\pipeline/md/b [54]), .ip3(n21335), 
        .ip4(n21334), .op(n8400) );
  nand2_1 U24141 ( .ip1(n21360), .ip2(n21336), .op(n21339) );
  nor2_1 U24142 ( .ip1(n21683), .ip2(n21336), .op(n21337) );
  nor2_1 U24143 ( .ip1(n21400), .ip2(n21337), .op(n21338) );
  mux2_1 U24144 ( .ip1(n21339), .ip2(n21338), .s(n22085), .op(n21342) );
  nand2_1 U24145 ( .ip1(\pipeline/md/b [51]), .ip2(n21493), .op(n21341) );
  nand2_1 U24146 ( .ip1(\pipeline/md/b [52]), .ip2(n14765), .op(n21340) );
  nand3_1 U24147 ( .ip1(n21342), .ip2(n21341), .ip3(n21340), .op(n8398) );
  nor2_1 U24148 ( .ip1(n21343), .ip2(n21414), .op(n21344) );
  xor2_1 U24149 ( .ip1(n21344), .ip2(n22084), .op(n21348) );
  nor2_1 U24150 ( .ip1(n21345), .ip2(n22665), .op(n21347) );
  nor2_1 U24151 ( .ip1(n22650), .ip2(n21680), .op(n21346) );
  ab_or_c_or_d U24152 ( .ip1(n22042), .ip2(n21348), .ip3(n21347), .ip4(n21346), 
        .op(n8395) );
  nand2_1 U24153 ( .ip1(n21427), .ip2(n21349), .op(n21350) );
  xor2_1 U24154 ( .ip1(n22083), .ip2(n21350), .op(n21351) );
  nor2_1 U24155 ( .ip1(n21351), .ip2(n21683), .op(n21353) );
  nor2_1 U24156 ( .ip1(n22650), .ip2(n22665), .op(n21352) );
  ab_or_c_or_d U24157 ( .ip1(n21493), .ip2(\pipeline/md/b [49]), .ip3(n21353), 
        .ip4(n21352), .op(n8394) );
  nor2_1 U24158 ( .ip1(n21354), .ip2(n21414), .op(n21355) );
  xor2_1 U24159 ( .ip1(n21355), .ip2(n17387), .op(n21356) );
  nand2_1 U24160 ( .ip1(n22042), .ip2(n21356), .op(n21359) );
  nand2_1 U24161 ( .ip1(\pipeline/md/b [49]), .ip2(n21440), .op(n21358) );
  nand2_1 U24162 ( .ip1(\pipeline/md/b [48]), .ip2(n21496), .op(n21357) );
  nand3_1 U24163 ( .ip1(n21359), .ip2(n21358), .ip3(n21357), .op(n8393) );
  nand2_1 U24164 ( .ip1(n21360), .ip2(n21361), .op(n21364) );
  nor2_1 U24165 ( .ip1(n21683), .ip2(n21361), .op(n21362) );
  nor2_1 U24166 ( .ip1(n21400), .ip2(n21362), .op(n21363) );
  mux2_1 U24167 ( .ip1(n21364), .ip2(n21363), .s(n22082), .op(n21367) );
  nand2_1 U24168 ( .ip1(\pipeline/md/b [47]), .ip2(n21493), .op(n21366) );
  nand2_1 U24169 ( .ip1(\pipeline/md/b [48]), .ip2(n14765), .op(n21365) );
  nand3_1 U24170 ( .ip1(n21367), .ip2(n21366), .ip3(n21365), .op(n8392) );
  nor2_1 U24171 ( .ip1(n22062), .ip2(n21374), .op(n21368) );
  nor2_1 U24172 ( .ip1(n21368), .ip2(n21414), .op(n21369) );
  xor2_1 U24173 ( .ip1(n21369), .ip2(n22064), .op(n21370) );
  nand2_1 U24174 ( .ip1(n22042), .ip2(n21370), .op(n21373) );
  nand2_1 U24175 ( .ip1(\pipeline/md/b [46]), .ip2(n21440), .op(n21372) );
  nand2_1 U24176 ( .ip1(\pipeline/md/b [45]), .ip2(n21496), .op(n21371) );
  nand3_1 U24177 ( .ip1(n21373), .ip2(n21372), .ip3(n21371), .op(n8387) );
  inv_1 U24178 ( .ip(n22062), .op(n21376) );
  nand2_1 U24179 ( .ip1(n21427), .ip2(n21374), .op(n21375) );
  xor2_1 U24180 ( .ip1(n21376), .ip2(n21375), .op(n21377) );
  nand2_1 U24181 ( .ip1(n22042), .ip2(n21377), .op(n21380) );
  nand2_1 U24182 ( .ip1(\pipeline/md/b [45]), .ip2(n20310), .op(n21379) );
  nand2_1 U24183 ( .ip1(\pipeline/md/b [44]), .ip2(n21493), .op(n21378) );
  nand3_1 U24184 ( .ip1(n21380), .ip2(n21379), .ip3(n21378), .op(n8386) );
  nor2_1 U24185 ( .ip1(n21381), .ip2(n21414), .op(n21382) );
  xor2_1 U24186 ( .ip1(n21383), .ip2(n21382), .op(n21384) );
  nor2_1 U24187 ( .ip1(n21384), .ip2(n21683), .op(n21386) );
  nor2_1 U24188 ( .ip1(n21390), .ip2(n21680), .op(n21385) );
  ab_or_c_or_d U24189 ( .ip1(n14765), .ip2(\pipeline/md/b [44]), .ip3(n21386), 
        .ip4(n21385), .op(n8385) );
  nand2_1 U24190 ( .ip1(n21427), .ip2(n21387), .op(n21388) );
  xor2_1 U24191 ( .ip1(n22058), .ip2(n21388), .op(n21389) );
  nor2_1 U24192 ( .ip1(n21389), .ip2(n21683), .op(n21392) );
  nor2_1 U24193 ( .ip1(n21390), .ip2(n22665), .op(n21391) );
  ab_or_c_or_d U24194 ( .ip1(n21493), .ip2(\pipeline/md/b [42]), .ip3(n21392), 
        .ip4(n21391), .op(n8384) );
  inv_1 U24195 ( .ip(n21393), .op(n21403) );
  nor2_1 U24196 ( .ip1(n21403), .ip2(n21406), .op(n21396) );
  nand2_1 U24197 ( .ip1(n22042), .ip2(n21403), .op(n21394) );
  nand2_1 U24198 ( .ip1(n21409), .ip2(n21394), .op(n21395) );
  mux2_1 U24199 ( .ip1(n21396), .ip2(n21395), .s(n22054), .op(n21398) );
  nor2_1 U24200 ( .ip1(n21763), .ip2(n22665), .op(n21397) );
  ab_or_c_or_d U24201 ( .ip1(n21493), .ip2(\pipeline/md/b [40]), .ip3(n21398), 
        .ip4(n21397), .op(n8377) );
  nand2_1 U24202 ( .ip1(n22042), .ip2(n21407), .op(n21408) );
  nor2_1 U24203 ( .ip1(n17376), .ip2(n21408), .op(n21399) );
  nor2_1 U24204 ( .ip1(n21400), .ip2(n21399), .op(n21401) );
  mux2_1 U24205 ( .ip1(n21406), .ip2(n21401), .s(n22052), .op(n21402) );
  nor2_1 U24206 ( .ip1(n21403), .ip2(n21402), .op(n21405) );
  nor2_1 U24207 ( .ip1(n21758), .ip2(n22665), .op(n21404) );
  ab_or_c_or_d U24208 ( .ip1(n21493), .ip2(\pipeline/md/b [39]), .ip3(n21405), 
        .ip4(n21404), .op(n8376) );
  nor2_1 U24209 ( .ip1(n21407), .ip2(n21406), .op(n21411) );
  nand2_1 U24210 ( .ip1(n21409), .ip2(n21408), .op(n21410) );
  mux2_1 U24211 ( .ip1(n21411), .ip2(n21410), .s(n17376), .op(n21413) );
  inv_1 U24212 ( .ip(\pipeline/md/b [38]), .op(n22553) );
  nor2_1 U24213 ( .ip1(n22553), .ip2(n21680), .op(n21412) );
  ab_or_c_or_d U24214 ( .ip1(n14765), .ip2(\pipeline/md/b [39]), .ip3(n21413), 
        .ip4(n21412), .op(n8374) );
  nor2_1 U24215 ( .ip1(n17370), .ip2(n21420), .op(n21415) );
  nor2_1 U24216 ( .ip1(n21415), .ip2(n21414), .op(n21416) );
  xor2_1 U24217 ( .ip1(n21416), .ip2(n22065), .op(n21419) );
  nor2_1 U24218 ( .ip1(n22553), .ip2(n22665), .op(n21418) );
  inv_1 U24219 ( .ip(\pipeline/md/b [37]), .op(n22543) );
  nor2_1 U24220 ( .ip1(n22543), .ip2(n21680), .op(n21417) );
  ab_or_c_or_d U24221 ( .ip1(n22042), .ip2(n21419), .ip3(n21418), .ip4(n21417), 
        .op(n8372) );
  nand2_1 U24222 ( .ip1(n21427), .ip2(n21420), .op(n21421) );
  xor2_1 U24223 ( .ip1(n17370), .ip2(n21421), .op(n21422) );
  nor2_1 U24224 ( .ip1(n21422), .ip2(n21683), .op(n21424) );
  nor2_1 U24225 ( .ip1(n22543), .ip2(n22665), .op(n21423) );
  ab_or_c_or_d U24226 ( .ip1(n21493), .ip2(\pipeline/md/b [36]), .ip3(n21424), 
        .ip4(n21423), .op(n8371) );
  nor2_1 U24227 ( .ip1(n22665), .ip2(n21425), .op(n21431) );
  nand2_1 U24228 ( .ip1(n21427), .ip2(n21426), .op(n21428) );
  xor2_1 U24229 ( .ip1(n22059), .ip2(n21428), .op(n21429) );
  nor2_1 U24230 ( .ip1(n21429), .ip2(n21683), .op(n21430) );
  ab_or_c_or_d U24231 ( .ip1(\pipeline/md/b [34]), .ip2(n21496), .ip3(n21431), 
        .ip4(n21430), .op(n8369) );
  nor2_1 U24232 ( .ip1(n22665), .ip2(n22484), .op(n21433) );
  nor2_1 U24233 ( .ip1(n21680), .ip2(n21656), .op(n21432) );
  ab_or_c_or_d U24234 ( .ip1(n22042), .ip2(n22053), .ip3(n21433), .ip4(n21432), 
        .op(n8365) );
  nand2_1 U24235 ( .ip1(n21440), .ip2(\pipeline/md/b [31]), .op(n21435) );
  nand2_1 U24236 ( .ip1(\pipeline/md/b [30]), .ip2(n21496), .op(n21434) );
  nand2_1 U24237 ( .ip1(n21435), .ip2(n21434), .op(n8364) );
  nand2_1 U24238 ( .ip1(n21440), .ip2(\pipeline/md/b [30]), .op(n21437) );
  nand2_1 U24239 ( .ip1(\pipeline/md/b [29]), .ip2(n21493), .op(n21436) );
  nand2_1 U24240 ( .ip1(n21437), .ip2(n21436), .op(n8363) );
  nand2_1 U24241 ( .ip1(n21440), .ip2(\pipeline/md/b [29]), .op(n21439) );
  nand2_1 U24242 ( .ip1(\pipeline/md/b [28]), .ip2(n21496), .op(n21438) );
  nand2_1 U24243 ( .ip1(n21439), .ip2(n21438), .op(n8362) );
  nand2_1 U24244 ( .ip1(n21440), .ip2(\pipeline/md/b [28]), .op(n21442) );
  nand2_1 U24245 ( .ip1(\pipeline/md/b [27]), .ip2(n21496), .op(n21441) );
  nand2_1 U24246 ( .ip1(n21442), .ip2(n21441), .op(n8361) );
  nand2_1 U24247 ( .ip1(n21440), .ip2(\pipeline/md/b [27]), .op(n21444) );
  nand2_1 U24248 ( .ip1(\pipeline/md/b [26]), .ip2(n21493), .op(n21443) );
  nand2_1 U24249 ( .ip1(n21444), .ip2(n21443), .op(n8360) );
  nand2_1 U24250 ( .ip1(n20310), .ip2(\pipeline/md/b [26]), .op(n21446) );
  nand2_1 U24251 ( .ip1(\pipeline/md/b [25]), .ip2(n21496), .op(n21445) );
  nand2_1 U24252 ( .ip1(n21446), .ip2(n21445), .op(n8359) );
  nand2_1 U24253 ( .ip1(n14765), .ip2(\pipeline/md/b [25]), .op(n21448) );
  nand2_1 U24254 ( .ip1(\pipeline/md/b [24]), .ip2(n21496), .op(n21447) );
  nand2_1 U24255 ( .ip1(n21448), .ip2(n21447), .op(n8358) );
  nand2_1 U24256 ( .ip1(n20310), .ip2(\pipeline/md/b [24]), .op(n21450) );
  nand2_1 U24257 ( .ip1(\pipeline/md/b [23]), .ip2(n21496), .op(n21449) );
  nand2_1 U24258 ( .ip1(n21450), .ip2(n21449), .op(n8357) );
  nand2_1 U24259 ( .ip1(n21440), .ip2(\pipeline/md/b [23]), .op(n21452) );
  nand2_1 U24260 ( .ip1(\pipeline/md/b [22]), .ip2(n21493), .op(n21451) );
  nand2_1 U24261 ( .ip1(n21452), .ip2(n21451), .op(n8356) );
  nand2_1 U24262 ( .ip1(n20310), .ip2(\pipeline/md/b [22]), .op(n21454) );
  nand2_1 U24263 ( .ip1(n21493), .ip2(\pipeline/md/b [21]), .op(n21453) );
  nand2_1 U24264 ( .ip1(n21454), .ip2(n21453), .op(n8355) );
  nand2_1 U24265 ( .ip1(n20310), .ip2(\pipeline/md/b [21]), .op(n21456) );
  nand2_1 U24266 ( .ip1(n21496), .ip2(\pipeline/md/b [20]), .op(n21455) );
  nand2_1 U24267 ( .ip1(n21456), .ip2(n21455), .op(n8354) );
  nand2_1 U24268 ( .ip1(n14765), .ip2(\pipeline/md/b [20]), .op(n21458) );
  nand2_1 U24269 ( .ip1(n21496), .ip2(\pipeline/md/b [19]), .op(n21457) );
  nand2_1 U24270 ( .ip1(n21458), .ip2(n21457), .op(n8353) );
  nand2_1 U24271 ( .ip1(n14765), .ip2(\pipeline/md/b [19]), .op(n21460) );
  nand2_1 U24272 ( .ip1(n21493), .ip2(\pipeline/md/b [18]), .op(n21459) );
  nand2_1 U24273 ( .ip1(n21460), .ip2(n21459), .op(n8352) );
  nand2_1 U24274 ( .ip1(n21440), .ip2(\pipeline/md/b [18]), .op(n21462) );
  nand2_1 U24275 ( .ip1(n21496), .ip2(\pipeline/md/b [17]), .op(n21461) );
  nand2_1 U24276 ( .ip1(n21462), .ip2(n21461), .op(n8351) );
  nand2_1 U24277 ( .ip1(n20310), .ip2(\pipeline/md/b [17]), .op(n21464) );
  nand2_1 U24278 ( .ip1(n21496), .ip2(\pipeline/md/b [16]), .op(n21463) );
  nand2_1 U24279 ( .ip1(n21464), .ip2(n21463), .op(n8350) );
  nand2_1 U24280 ( .ip1(n14765), .ip2(\pipeline/md/b [16]), .op(n21466) );
  nand2_1 U24281 ( .ip1(n21496), .ip2(\pipeline/md/b [15]), .op(n21465) );
  nand2_1 U24282 ( .ip1(n21466), .ip2(n21465), .op(n8349) );
  nand2_1 U24283 ( .ip1(n20310), .ip2(\pipeline/md/b [15]), .op(n21468) );
  nand2_1 U24284 ( .ip1(n21493), .ip2(\pipeline/md/b [14]), .op(n21467) );
  nand2_1 U24285 ( .ip1(n21468), .ip2(n21467), .op(n8348) );
  nand2_1 U24286 ( .ip1(n14765), .ip2(\pipeline/md/b [14]), .op(n21470) );
  nand2_1 U24287 ( .ip1(n21496), .ip2(\pipeline/md/b [13]), .op(n21469) );
  nand2_1 U24288 ( .ip1(n21470), .ip2(n21469), .op(n8347) );
  nand2_1 U24289 ( .ip1(n21440), .ip2(\pipeline/md/b [13]), .op(n21472) );
  nand2_1 U24290 ( .ip1(n21496), .ip2(\pipeline/md/b [12]), .op(n21471) );
  nand2_1 U24291 ( .ip1(n21472), .ip2(n21471), .op(n8346) );
  nand2_1 U24292 ( .ip1(n14765), .ip2(\pipeline/md/b [12]), .op(n21474) );
  nand2_1 U24293 ( .ip1(n21493), .ip2(\pipeline/md/b [11]), .op(n21473) );
  nand2_1 U24294 ( .ip1(n21474), .ip2(n21473), .op(n8345) );
  nand2_1 U24295 ( .ip1(n20310), .ip2(\pipeline/md/b [11]), .op(n21476) );
  nand2_1 U24296 ( .ip1(n21496), .ip2(\pipeline/md/b [10]), .op(n21475) );
  nand2_1 U24297 ( .ip1(n21476), .ip2(n21475), .op(n8344) );
  nand2_1 U24298 ( .ip1(n14765), .ip2(\pipeline/md/b [10]), .op(n21478) );
  nand2_1 U24299 ( .ip1(n21496), .ip2(\pipeline/md/b [9]), .op(n21477) );
  nand2_1 U24300 ( .ip1(n21478), .ip2(n21477), .op(n8343) );
  nand2_1 U24301 ( .ip1(n21440), .ip2(\pipeline/md/b [9]), .op(n21480) );
  nand2_1 U24302 ( .ip1(n21496), .ip2(\pipeline/md/b [8]), .op(n21479) );
  nand2_1 U24303 ( .ip1(n21480), .ip2(n21479), .op(n8342) );
  nand2_1 U24304 ( .ip1(n20310), .ip2(\pipeline/md/b [8]), .op(n21482) );
  nand2_1 U24305 ( .ip1(n21493), .ip2(\pipeline/md/b [7]), .op(n21481) );
  nand2_1 U24306 ( .ip1(n21482), .ip2(n21481), .op(n8341) );
  nand2_1 U24307 ( .ip1(n14765), .ip2(\pipeline/md/b [7]), .op(n21484) );
  nand2_1 U24308 ( .ip1(n21496), .ip2(\pipeline/md/b [6]), .op(n21483) );
  nand2_1 U24309 ( .ip1(n21484), .ip2(n21483), .op(n8340) );
  nand2_1 U24310 ( .ip1(n21440), .ip2(\pipeline/md/b [6]), .op(n21486) );
  nand2_1 U24311 ( .ip1(n21496), .ip2(\pipeline/md/b [5]), .op(n21485) );
  nand2_1 U24312 ( .ip1(n21486), .ip2(n21485), .op(n8339) );
  nand2_1 U24313 ( .ip1(n20310), .ip2(\pipeline/md/b [5]), .op(n21488) );
  nand2_1 U24314 ( .ip1(n21493), .ip2(\pipeline/md/b [4]), .op(n21487) );
  nand2_1 U24315 ( .ip1(n21488), .ip2(n21487), .op(n8338) );
  nand2_1 U24316 ( .ip1(n14765), .ip2(\pipeline/md/b [4]), .op(n21490) );
  nand2_1 U24317 ( .ip1(n21493), .ip2(\pipeline/md/b [3]), .op(n21489) );
  nand2_1 U24318 ( .ip1(n21490), .ip2(n21489), .op(n8337) );
  nand2_1 U24319 ( .ip1(n21440), .ip2(\pipeline/md/b [3]), .op(n21492) );
  nand2_1 U24320 ( .ip1(n21496), .ip2(\pipeline/md/b [2]), .op(n21491) );
  nand2_1 U24321 ( .ip1(n21492), .ip2(n21491), .op(n8336) );
  nand2_1 U24322 ( .ip1(n21440), .ip2(\pipeline/md/b [2]), .op(n21495) );
  nand2_1 U24323 ( .ip1(n21493), .ip2(\pipeline/md/b [1]), .op(n21494) );
  nand2_1 U24324 ( .ip1(n21495), .ip2(n21494), .op(n8335) );
  nand2_1 U24325 ( .ip1(n14765), .ip2(\pipeline/md/b [1]), .op(n21498) );
  nand2_1 U24326 ( .ip1(n21496), .ip2(\pipeline/md/b [0]), .op(n21497) );
  nand2_1 U24327 ( .ip1(n21498), .ip2(n21497), .op(n8334) );
  or2_1 U24328 ( .ip1(\pipeline/md/b [0]), .ip2(n22665), .op(n21521) );
  nand2_1 U24329 ( .ip1(n14770), .ip2(n21521), .op(n21504) );
  nor2_1 U24330 ( .ip1(n21500), .ip2(n21499), .op(n21503) );
  nor2_1 U24331 ( .ip1(n21730), .ip2(n21501), .op(n21502) );
  ab_or_c_or_d U24332 ( .ip1(\pipeline/md/a [0]), .ip2(n21504), .ip3(n21503), 
        .ip4(n21502), .op(n8426) );
  nor3_1 U24333 ( .ip1(\pipeline/md/result [32]), .ip2(n21506), .ip3(n21505), 
        .op(n21513) );
  inv_1 U24334 ( .ip(n21506), .op(n21507) );
  nor2_1 U24335 ( .ip1(n21662), .ip2(n21507), .op(n21508) );
  nor2_1 U24336 ( .ip1(n21509), .ip2(n21508), .op(n21511) );
  nor2_1 U24337 ( .ip1(n21511), .ip2(n21510), .op(n21512) );
  nor2_1 U24338 ( .ip1(n21513), .ip2(n21512), .op(n21514) );
  nor2_1 U24339 ( .ip1(n21514), .ip2(n21967), .op(n21519) );
  nor3_1 U24340 ( .ip1(n21517), .ip2(n21516), .ip3(n21515), .op(n21518) );
  not_ab_or_c_or_d U24341 ( .ip1(n21972), .ip2(n21520), .ip3(n21519), .ip4(
        n21518), .op(n21526) );
  nand2_1 U24342 ( .ip1(n22738), .ip2(n21521), .op(n21522) );
  nand2_1 U24343 ( .ip1(\pipeline/md_resp_result [0]), .ip2(n21522), .op(
        n21525) );
  nand3_1 U24344 ( .ip1(n22750), .ip2(\pipeline/md/b [0]), .ip3(n21523), .op(
        n21524) );
  nand3_1 U24345 ( .ip1(n21526), .ip2(n21525), .ip3(n21524), .op(n8634) );
  mux2_1 U24346 ( .ip1(\pipeline/csr_rdata_WB [0]), .ip2(n21527), .s(n17429), 
        .op(n8806) );
  inv_1 U24347 ( .ip(n21528), .op(n21529) );
  nand3_1 U24348 ( .ip1(n21531), .ip2(n21530), .ip3(n21529), .op(n21581) );
  nand2_1 U24349 ( .ip1(n21533), .ip2(n21532), .op(n21535) );
  nand2_1 U24350 ( .ip1(n21535), .ip2(n21534), .op(n21539) );
  nand2_1 U24351 ( .ip1(n21536), .ip2(n13728), .op(n21538) );
  nand2_1 U24352 ( .ip1(n21541), .ip2(n21540), .op(n21542) );
  nand2_1 U24353 ( .ip1(n21543), .ip2(n21542), .op(n21571) );
  nand2_1 U24354 ( .ip1(n21544), .ip2(n16776), .op(n21546) );
  nor4_1 U24355 ( .ip1(n21548), .ip2(n21547), .ip3(n21546), .ip4(n21545), .op(
        n21570) );
  nand2_1 U24356 ( .ip1(n21550), .ip2(n21549), .op(n21568) );
  nor3_1 U24357 ( .ip1(n21553), .ip2(n21551), .ip3(n13870), .op(n21561) );
  nor2_1 U24358 ( .ip1(n21552), .ip2(n13524), .op(n21559) );
  nor2_1 U24359 ( .ip1(n21553), .ip2(n13870), .op(n21554) );
  nor2_1 U24360 ( .ip1(n21555), .ip2(n21554), .op(n21556) );
  nor2_1 U24361 ( .ip1(n21557), .ip2(n21556), .op(n21558) );
  nor2_1 U24362 ( .ip1(n21559), .ip2(n21558), .op(n21560) );
  not_ab_or_c_or_d U24363 ( .ip1(n21563), .ip2(n21562), .ip3(n21561), .ip4(
        n21560), .op(n21567) );
  or2_1 U24364 ( .ip1(n21565), .ip2(n21564), .op(n21566) );
  nand3_1 U24365 ( .ip1(n21568), .ip2(n21567), .ip3(n21566), .op(n21569) );
  not_ab_or_c_or_d U24366 ( .ip1(n21572), .ip2(n21571), .ip3(n21570), .ip4(
        n21569), .op(n21580) );
  nand2_1 U24367 ( .ip1(n21574), .ip2(n21573), .op(n21576) );
  xnor2_1 U24368 ( .ip1(n21576), .ip2(n21575), .op(n21578) );
  nand2_1 U24369 ( .ip1(n21578), .ip2(n21577), .op(n21579) );
  nand3_1 U24370 ( .ip1(n21581), .ip2(n21580), .ip3(n21579), .op(dmem_haddr[0]) );
  mux2_1 U24371 ( .ip1(dmem_haddr[0]), .ip2(\pipeline/alu_out_WB [0]), .s(
        n21582), .op(n8807) );
  nand2_1 U24372 ( .ip1(n21584), .ip2(n21583), .op(n21587) );
  nand2_1 U24373 ( .ip1(dmem_rdata[31]), .ip2(n21585), .op(n21586) );
  nand3_1 U24374 ( .ip1(n21588), .ip2(n21587), .ip3(n21586), .op(n21620) );
  mux2_1 U24375 ( .ip1(\pipeline/regfile/data[22][31] ), .ip2(n21620), .s(
        n21589), .op(n9193) );
  mux2_1 U24376 ( .ip1(\pipeline/regfile/data[28][31] ), .ip2(n21620), .s(
        n21590), .op(n9001) );
  mux2_1 U24377 ( .ip1(\pipeline/regfile/data[12][31] ), .ip2(n21620), .s(
        n21591), .op(n9513) );
  mux2_1 U24378 ( .ip1(\pipeline/regfile/data[19][31] ), .ip2(n21620), .s(
        n21592), .op(n9289) );
  mux2_1 U24379 ( .ip1(\pipeline/regfile/data[11][31] ), .ip2(n21620), .s(
        n21593), .op(n9545) );
  mux2_1 U24380 ( .ip1(\pipeline/regfile/data[30][31] ), .ip2(n21620), .s(
        n21594), .op(n8937) );
  mux2_1 U24381 ( .ip1(\pipeline/regfile/data[18][31] ), .ip2(n21620), .s(
        n21595), .op(n9321) );
  mux2_1 U24382 ( .ip1(\pipeline/regfile/data[23][31] ), .ip2(n21620), .s(
        n21596), .op(n9161) );
  mux2_1 U24383 ( .ip1(\pipeline/regfile/data[6][31] ), .ip2(n21620), .s(
        n21597), .op(n9705) );
  mux2_1 U24384 ( .ip1(\pipeline/regfile/data[5][31] ), .ip2(n21620), .s(
        n21598), .op(n9737) );
  mux2_1 U24385 ( .ip1(\pipeline/regfile/data[3][31] ), .ip2(n21620), .s(
        n21599), .op(n9801) );
  mux2_1 U24386 ( .ip1(\pipeline/regfile/data[13][31] ), .ip2(n21620), .s(
        n21600), .op(n9481) );
  mux2_1 U24387 ( .ip1(\pipeline/regfile/data[20][31] ), .ip2(n21620), .s(
        n21601), .op(n9257) );
  mux2_1 U24388 ( .ip1(\pipeline/regfile/data[25][31] ), .ip2(n21620), .s(
        n21602), .op(n9097) );
  mux2_1 U24389 ( .ip1(\pipeline/regfile/data[24][31] ), .ip2(n21620), .s(
        n21603), .op(n9129) );
  mux2_1 U24390 ( .ip1(\pipeline/regfile/data[14][31] ), .ip2(n21620), .s(
        n21604), .op(n9449) );
  mux2_1 U24391 ( .ip1(\pipeline/regfile/data[4][31] ), .ip2(n21620), .s(
        n21605), .op(n9769) );
  mux2_1 U24392 ( .ip1(\pipeline/regfile/data[31][31] ), .ip2(n21620), .s(
        n21606), .op(n8905) );
  mux2_1 U24393 ( .ip1(\pipeline/regfile/data[26][31] ), .ip2(n21620), .s(
        n21607), .op(n9065) );
  mux2_1 U24394 ( .ip1(\pipeline/regfile/data[16][31] ), .ip2(n21620), .s(
        n21608), .op(n9385) );
  mux2_1 U24395 ( .ip1(\pipeline/regfile/data[9][31] ), .ip2(n21620), .s(
        n21609), .op(n9609) );
  mux2_1 U24396 ( .ip1(\pipeline/regfile/data[2][31] ), .ip2(n21620), .s(
        n21610), .op(n9833) );
  mux2_1 U24397 ( .ip1(\pipeline/regfile/data[1][31] ), .ip2(n21620), .s(
        n21611), .op(n9865) );
  mux2_1 U24398 ( .ip1(\pipeline/regfile/data[27][31] ), .ip2(n21620), .s(
        n21612), .op(n9033) );
  mux2_1 U24399 ( .ip1(\pipeline/regfile/data[15][31] ), .ip2(n21620), .s(
        n21613), .op(n9417) );
  mux2_1 U24400 ( .ip1(\pipeline/regfile/data[7][31] ), .ip2(n21620), .s(
        n21614), .op(n9673) );
  mux2_1 U24401 ( .ip1(\pipeline/regfile/data[21][31] ), .ip2(n21620), .s(
        n21615), .op(n9225) );
  mux2_1 U24402 ( .ip1(\pipeline/regfile/data[17][31] ), .ip2(n21620), .s(
        n21616), .op(n9353) );
  mux2_1 U24403 ( .ip1(\pipeline/regfile/data[8][31] ), .ip2(n21620), .s(
        n21617), .op(n9641) );
  mux2_1 U24404 ( .ip1(\pipeline/regfile/data[10][31] ), .ip2(n21620), .s(
        n21618), .op(n9577) );
  mux2_1 U24405 ( .ip1(\pipeline/regfile/data[29][31] ), .ip2(n21620), .s(
        n21619), .op(n8969) );
  nand2_1 U24406 ( .ip1(n21622), .ip2(n21621), .op(n21623) );
  nand2_1 U24407 ( .ip1(n21624), .ip2(n21623), .op(n21648) );
  xor2_1 U24408 ( .ip1(n21625), .ip2(n21648), .op(n21626) );
  nand2_1 U24409 ( .ip1(n21649), .ip2(n21626), .op(n21635) );
  nand2_1 U24410 ( .ip1(n21628), .ip2(n21627), .op(n21629) );
  nand2_1 U24411 ( .ip1(n21630), .ip2(n21629), .op(n21636) );
  xor2_1 U24412 ( .ip1(\pipeline/md/b [30]), .ip2(n21636), .op(n21631) );
  nor2_1 U24413 ( .ip1(n21947), .ip2(n21631), .op(n21632) );
  xor2_1 U24414 ( .ip1(\pipeline/md/a [30]), .ip2(n21632), .op(n21633) );
  nand2_1 U24415 ( .ip1(n21633), .ip2(n21643), .op(n21634) );
  nand2_1 U24416 ( .ip1(n21635), .ip2(n21634), .op(n8421) );
  inv_1 U24417 ( .ip(n21636), .op(n21638) );
  nor2_1 U24418 ( .ip1(n21638), .ip2(n21637), .op(n21695) );
  nor2_1 U24419 ( .ip1(n21695), .ip2(n21639), .op(n21640) );
  xor2_1 U24420 ( .ip1(n21640), .ip2(n21656), .op(n21641) );
  nor2_1 U24421 ( .ip1(n21947), .ip2(n21641), .op(n21642) );
  xor2_1 U24422 ( .ip1(\pipeline/md/a [31]), .ip2(n21642), .op(n21644) );
  nand2_1 U24423 ( .ip1(n21644), .ip2(n21643), .op(n21651) );
  nand2_1 U24424 ( .ip1(n21646), .ip2(n21645), .op(n21647) );
  nand4_1 U24425 ( .ip1(n21649), .ip2(n14594), .ip3(n21648), .ip4(n21647), 
        .op(n21650) );
  nand2_1 U24426 ( .ip1(n21651), .ip2(n21650), .op(n8521) );
  nor2_1 U24427 ( .ip1(\pipeline/md_resp_result [30]), .ip2(n21652), .op(
        n21653) );
  or2_1 U24428 ( .ip1(n21654), .ip2(n21653), .op(n21657) );
  inv_1 U24429 ( .ip(n21657), .op(n21655) );
  nor2_1 U24430 ( .ip1(\pipeline/md/b [31]), .ip2(n21655), .op(n22485) );
  nor2_1 U24431 ( .ip1(n21657), .ip2(n21656), .op(n22482) );
  nor4_1 U24432 ( .ip1(\pipeline/md_resp_result [31]), .ip2(n22485), .ip3(
        n22482), .ip4(n22755), .op(n21670) );
  nor2_1 U24433 ( .ip1(n21658), .ip2(n21957), .op(n21667) );
  nor3_1 U24434 ( .ip1(n21666), .ip2(n21960), .ip3(n21667), .op(n21665) );
  nor2_1 U24435 ( .ip1(n21660), .ip2(n21659), .op(n21663) );
  nor2_1 U24436 ( .ip1(\pipeline/md/result [63]), .ip2(n21663), .op(n21661) );
  not_ab_or_c_or_d U24437 ( .ip1(\pipeline/md/result [63]), .ip2(n21663), 
        .ip3(n21662), .ip4(n21661), .op(n21664) );
  not_ab_or_c_or_d U24438 ( .ip1(n21667), .ip2(n21666), .ip3(n21665), .ip4(
        n21664), .op(n21668) );
  nor2_1 U24439 ( .ip1(n21668), .ip2(n21967), .op(n21669) );
  not_ab_or_c_or_d U24440 ( .ip1(n21672), .ip2(n21671), .ip3(n21670), .ip4(
        n21669), .op(n21677) );
  or2_1 U24441 ( .ip1(n22485), .ip2(n22482), .op(n21673) );
  nand2_1 U24442 ( .ip1(n20310), .ip2(n21673), .op(n21674) );
  nand2_1 U24443 ( .ip1(n22738), .ip2(n21674), .op(n21675) );
  nand2_1 U24444 ( .ip1(\pipeline/md_resp_result [31]), .ip2(n21675), .op(
        n21676) );
  nand2_1 U24445 ( .ip1(n21677), .ip2(n21676), .op(n8603) );
  inv_1 U24446 ( .ip(n21678), .op(n21679) );
  mux2_1 U24447 ( .ip1(\pipeline/csr_rdata_WB [31]), .ip2(n21679), .s(n17429), 
        .op(n10072) );
  nor2_1 U24448 ( .ip1(n21681), .ip2(n21680), .op(n21688) );
  inv_1 U24449 ( .ip(n21682), .op(n21685) );
  inv_1 U24450 ( .ip(n22069), .op(n21684) );
  not_ab_or_c_or_d U24451 ( .ip1(n21686), .ip2(n21685), .ip3(n21684), .ip4(
        n21683), .op(n21687) );
  or2_1 U24452 ( .ip1(n21688), .ip2(n21687), .op(n8496) );
  nand2_1 U24453 ( .ip1(\pipeline/md/a [60]), .ip2(n21884), .op(n21733) );
  inv_1 U24454 ( .ip(n21885), .op(n21719) );
  inv_1 U24455 ( .ip(\pipeline/md/a [50]), .op(n21740) );
  inv_1 U24456 ( .ip(n21689), .op(n21713) );
  inv_1 U24457 ( .ip(n21690), .op(n21710) );
  inv_1 U24458 ( .ip(n21691), .op(n21704) );
  inv_1 U24459 ( .ip(n21692), .op(n21813) );
  inv_1 U24460 ( .ip(n21693), .op(n21699) );
  nor2_1 U24461 ( .ip1(n21695), .ip2(n21694), .op(n21696) );
  or2_1 U24462 ( .ip1(n21697), .ip2(n21696), .op(n21795) );
  nand3_1 U24463 ( .ip1(n21795), .ip2(n21794), .ip3(n21799), .op(n21698) );
  nand2_1 U24464 ( .ip1(n21699), .ip2(n21698), .op(n21772) );
  inv_1 U24465 ( .ip(n21808), .op(n21700) );
  nand2_1 U24466 ( .ip1(n21806), .ip2(n21700), .op(n21814) );
  and2_1 U24467 ( .ip1(n21701), .ip2(n21814), .op(n21702) );
  nor2_1 U24468 ( .ip1(n21813), .ip2(n21702), .op(n21757) );
  nor3_1 U24469 ( .ip1(n21704), .ip2(n21757), .ip3(n21703), .op(n21706) );
  nor2_1 U24470 ( .ip1(n21706), .ip2(n21705), .op(n21833) );
  nand2_1 U24471 ( .ip1(n21833), .ip2(n21831), .op(n21707) );
  nand2_1 U24472 ( .ip1(n21832), .ip2(n21707), .op(n21841) );
  nand2_1 U24473 ( .ip1(n21839), .ip2(n21841), .op(n21847) );
  nand2_1 U24474 ( .ip1(n21708), .ip2(n21847), .op(n21709) );
  nand2_1 U24475 ( .ip1(n21710), .ip2(n21709), .op(n21854) );
  nand2_1 U24476 ( .ip1(n21711), .ip2(n21854), .op(n21712) );
  nand2_1 U24477 ( .ip1(n21713), .ip2(n21712), .op(n21862) );
  nand2_1 U24478 ( .ip1(n21714), .ip2(n21862), .op(n21715) );
  nand2_1 U24479 ( .ip1(n21716), .ip2(n21715), .op(n21749) );
  nor2_1 U24480 ( .ip1(n21867), .ip2(n21870), .op(n21875) );
  or2_1 U24481 ( .ip1(n21875), .ip2(n21717), .op(n21718) );
  nand2_1 U24482 ( .ip1(n21877), .ip2(n21718), .op(n21887) );
  nor2_1 U24483 ( .ip1(n21719), .ip2(n21887), .op(n21892) );
  nor2_1 U24484 ( .ip1(n21892), .ip2(n21720), .op(n21721) );
  nor2_1 U24485 ( .ip1(n21894), .ip2(n21721), .op(n21909) );
  nor2_1 U24486 ( .ip1(n21909), .ip2(n21904), .op(n21722) );
  nor2_1 U24487 ( .ip1(n21723), .ip2(n21722), .op(n21917) );
  nor2_1 U24488 ( .ip1(n21917), .ip2(n21918), .op(n21724) );
  nor2_1 U24489 ( .ip1(n21725), .ip2(n21724), .op(n21937) );
  inv_1 U24490 ( .ip(n21937), .op(n21726) );
  nand3_1 U24491 ( .ip1(n21936), .ip2(n21727), .ip3(n21726), .op(n21728) );
  nand2_1 U24492 ( .ip1(n21729), .ip2(n21728), .op(n21734) );
  or2_1 U24493 ( .ip1(n21731), .ip2(n21730), .op(n21732) );
  nand2_1 U24494 ( .ip1(n21733), .ip2(n21732), .op(n8542) );
  nand2_1 U24495 ( .ip1(\pipeline/md/a [61]), .ip2(n21947), .op(n21738) );
  inv_1 U24496 ( .ip(\pipeline/md/a [61]), .op(n21949) );
  fulladder U24497 ( .a(\pipeline/md/b [60]), .b(n21735), .ci(n21734), .co(
        n21948), .s(n21731) );
  or2_1 U24498 ( .ip1(n21736), .ip2(n21730), .op(n21737) );
  nand2_1 U24499 ( .ip1(n21738), .ip2(n21737), .op(n8541) );
  nand2_1 U24500 ( .ip1(\pipeline/md/a [50]), .ip2(n21884), .op(n21743) );
  fulladder U24501 ( .a(\pipeline/md/b [50]), .b(n21740), .ci(n21739), .co(
        n21744), .s(n21741) );
  or2_1 U24502 ( .ip1(n21741), .ip2(n21730), .op(n21742) );
  nand2_1 U24503 ( .ip1(n21743), .ip2(n21742), .op(n8552) );
  nand2_1 U24504 ( .ip1(\pipeline/md/a [51]), .ip2(n21947), .op(n21748) );
  fulladder U24505 ( .a(n21745), .b(\pipeline/md/b [51]), .ci(n21744), .co(
        n21870), .s(n21746) );
  or2_1 U24506 ( .ip1(n21746), .ip2(n21730), .op(n21747) );
  nand2_1 U24507 ( .ip1(n21748), .ip2(n21747), .op(n8551) );
  nand2_1 U24508 ( .ip1(\pipeline/md/a [49]), .ip2(n21884), .op(n21753) );
  fulladder U24509 ( .a(n21750), .b(\pipeline/md/b [49]), .ci(n21749), .co(
        n21739), .s(n21751) );
  or2_1 U24510 ( .ip1(n21751), .ip2(n21730), .op(n21752) );
  nand2_1 U24511 ( .ip1(n21753), .ip2(n21752), .op(n8553) );
  nand2_1 U24512 ( .ip1(\pipeline/md/a [42]), .ip2(n21884), .op(n21756) );
  nand2_1 U24513 ( .ip1(n21944), .ip2(n21754), .op(n21755) );
  nand2_1 U24514 ( .ip1(n21756), .ip2(n21755), .op(n8560) );
  nand2_1 U24515 ( .ip1(\pipeline/md/a [40]), .ip2(n21947), .op(n21761) );
  fulladder U24516 ( .a(n21758), .b(\pipeline/md/a [40]), .ci(n21757), .co(
        n21762), .s(n21759) );
  nand2_1 U24517 ( .ip1(n21944), .ip2(n21759), .op(n21760) );
  nand2_1 U24518 ( .ip1(n21761), .ip2(n21760), .op(n8562) );
  nand2_1 U24519 ( .ip1(\pipeline/md/a [41]), .ip2(n21884), .op(n21766) );
  fulladder U24520 ( .a(\pipeline/md/a [41]), .b(n21763), .ci(n21762), .co(
        n21821), .s(n21764) );
  nand2_1 U24521 ( .ip1(n21944), .ip2(n21764), .op(n21765) );
  nand2_1 U24522 ( .ip1(n21766), .ip2(n21765), .op(n8561) );
  nand2_1 U24523 ( .ip1(n21947), .ip2(\pipeline/md/a [36]), .op(n21771) );
  fulladder U24524 ( .a(\pipeline/md/b [36]), .b(n21768), .ci(n21767), .co(
        n21777), .s(n21769) );
  or2_1 U24525 ( .ip1(n21769), .ip2(n21730), .op(n21770) );
  nand2_1 U24526 ( .ip1(n21771), .ip2(n21770), .op(n8566) );
  nand2_1 U24527 ( .ip1(n21884), .ip2(\pipeline/md/a [34]), .op(n21776) );
  fulladder U24528 ( .a(\pipeline/md/b [34]), .b(n21773), .ci(n21772), .co(
        n21782), .s(n21774) );
  or2_1 U24529 ( .ip1(n21774), .ip2(n21730), .op(n21775) );
  nand2_1 U24530 ( .ip1(n21776), .ip2(n21775), .op(n8568) );
  nand2_1 U24531 ( .ip1(\pipeline/md/a [37]), .ip2(n21884), .op(n21781) );
  fulladder U24532 ( .a(n21778), .b(\pipeline/md/b [37]), .ci(n21777), .co(
        n21808), .s(n21779) );
  or2_1 U24533 ( .ip1(n21779), .ip2(n21730), .op(n21780) );
  nand2_1 U24534 ( .ip1(n21781), .ip2(n21780), .op(n8565) );
  nand2_1 U24535 ( .ip1(n21947), .ip2(\pipeline/md/a [35]), .op(n21786) );
  fulladder U24536 ( .a(n21783), .b(\pipeline/md/b [35]), .ci(n21782), .co(
        n21767), .s(n21784) );
  or2_1 U24537 ( .ip1(n21784), .ip2(n21730), .op(n21785) );
  nand2_1 U24538 ( .ip1(n21786), .ip2(n21785), .op(n8567) );
  xor2_1 U24539 ( .ip1(\pipeline/md/b [32]), .ip2(n21795), .op(n21790) );
  inv_1 U24540 ( .ip(n21790), .op(n21787) );
  nand2_1 U24541 ( .ip1(n21440), .ip2(n21787), .op(n21788) );
  nand2_1 U24542 ( .ip1(n14770), .ip2(n21788), .op(n21789) );
  nand2_1 U24543 ( .ip1(\pipeline/md/a [32]), .ip2(n21789), .op(n21793) );
  nand3_1 U24544 ( .ip1(n21944), .ip2(n21791), .ip3(n21790), .op(n21792) );
  nand2_1 U24545 ( .ip1(n21793), .ip2(n21792), .op(n8570) );
  nand2_1 U24546 ( .ip1(n21884), .ip2(\pipeline/md/a [33]), .op(n21804) );
  nand2_1 U24547 ( .ip1(n21795), .ip2(n21794), .op(n21796) );
  nand2_1 U24548 ( .ip1(n21797), .ip2(n21796), .op(n21801) );
  nand2_1 U24549 ( .ip1(n21799), .ip2(n21798), .op(n21800) );
  xor2_1 U24550 ( .ip1(n21801), .ip2(n21800), .op(n21802) );
  nand2_1 U24551 ( .ip1(n21944), .ip2(n21802), .op(n21803) );
  nand2_1 U24552 ( .ip1(n21804), .ip2(n21803), .op(n8569) );
  nand2_1 U24553 ( .ip1(\pipeline/md/a [38]), .ip2(n21884), .op(n21811) );
  inv_1 U24554 ( .ip(n21805), .op(n21815) );
  nand2_1 U24555 ( .ip1(n21806), .ip2(n21815), .op(n21807) );
  xor2_1 U24556 ( .ip1(n21808), .ip2(n21807), .op(n21809) );
  nand2_1 U24557 ( .ip1(n21944), .ip2(n21809), .op(n21810) );
  nand2_1 U24558 ( .ip1(n21811), .ip2(n21810), .op(n8564) );
  nand2_1 U24559 ( .ip1(\pipeline/md/a [39]), .ip2(n21947), .op(n21820) );
  nor2_1 U24560 ( .ip1(n21813), .ip2(n21812), .op(n21817) );
  nand2_1 U24561 ( .ip1(n21815), .ip2(n21814), .op(n21816) );
  xor2_1 U24562 ( .ip1(n21817), .ip2(n21816), .op(n21818) );
  nand2_1 U24563 ( .ip1(n21944), .ip2(n21818), .op(n21819) );
  nand2_1 U24564 ( .ip1(n21820), .ip2(n21819), .op(n8563) );
  nand2_1 U24565 ( .ip1(\pipeline/md/a [43]), .ip2(n21884), .op(n21829) );
  fulladder U24566 ( .a(n21822), .b(\pipeline/md/a [42]), .ci(n21821), .co(
        n21826), .s(n21754) );
  nor2_1 U24567 ( .ip1(n21824), .ip2(n21823), .op(n21825) );
  xor2_1 U24568 ( .ip1(n21826), .ip2(n21825), .op(n21827) );
  nand2_1 U24569 ( .ip1(n21944), .ip2(n21827), .op(n21828) );
  nand2_1 U24570 ( .ip1(n21829), .ip2(n21828), .op(n8559) );
  nand2_1 U24571 ( .ip1(\pipeline/md/a [44]), .ip2(n21947), .op(n21838) );
  xor2_1 U24572 ( .ip1(\pipeline/md/b [44]), .ip2(n21830), .op(n21835) );
  nand2_1 U24573 ( .ip1(n21832), .ip2(n21831), .op(n21834) );
  mux2_1 U24574 ( .ip1(n21835), .ip2(n21834), .s(n21833), .op(n21836) );
  nand2_1 U24575 ( .ip1(n21944), .ip2(n21836), .op(n21837) );
  nand2_1 U24576 ( .ip1(n21838), .ip2(n21837), .op(n8558) );
  nand2_1 U24577 ( .ip1(\pipeline/md/a [45]), .ip2(n21947), .op(n21845) );
  inv_1 U24578 ( .ip(n21839), .op(n21840) );
  nor2_1 U24579 ( .ip1(n21840), .ip2(n21846), .op(n21842) );
  xor2_1 U24580 ( .ip1(n21842), .ip2(n21841), .op(n21843) );
  nand2_1 U24581 ( .ip1(n21944), .ip2(n21843), .op(n21844) );
  nand2_1 U24582 ( .ip1(n21845), .ip2(n21844), .op(n8557) );
  inv_1 U24583 ( .ip(n21846), .op(n21848) );
  nand2_1 U24584 ( .ip1(n21848), .ip2(n21847), .op(n21849) );
  xor2_1 U24585 ( .ip1(\pipeline/md/b [46]), .ip2(n21849), .op(n21850) );
  nor2_1 U24586 ( .ip1(n21884), .ip2(n21850), .op(n21852) );
  xor2_1 U24587 ( .ip1(n21852), .ip2(n21851), .op(n21853) );
  nor2_1 U24588 ( .ip1(n21866), .ip2(n21853), .op(n8556) );
  xor2_1 U24589 ( .ip1(\pipeline/md/b [47]), .ip2(n21854), .op(n21858) );
  inv_1 U24590 ( .ip(n21858), .op(n21855) );
  nand2_1 U24591 ( .ip1(n20310), .ip2(n21855), .op(n21856) );
  nand2_1 U24592 ( .ip1(n14770), .ip2(n21856), .op(n21857) );
  nand2_1 U24593 ( .ip1(\pipeline/md/a [47]), .ip2(n21857), .op(n21861) );
  inv_1 U24594 ( .ip(\pipeline/md/a [47]), .op(n21859) );
  nand3_1 U24595 ( .ip1(n21944), .ip2(n21859), .ip3(n21858), .op(n21860) );
  nand2_1 U24596 ( .ip1(n21861), .ip2(n21860), .op(n8555) );
  xor2_1 U24597 ( .ip1(\pipeline/md/b [48]), .ip2(n21862), .op(n21863) );
  nand2_1 U24598 ( .ip1(n14770), .ip2(n21863), .op(n21864) );
  xor2_1 U24599 ( .ip1(\pipeline/md/a [48]), .ip2(n21864), .op(n21865) );
  nor2_1 U24600 ( .ip1(n21866), .ip2(n21865), .op(n8554) );
  nand2_1 U24601 ( .ip1(\pipeline/md/a [52]), .ip2(n21947), .op(n21873) );
  inv_1 U24602 ( .ip(n21867), .op(n21868) );
  nand2_1 U24603 ( .ip1(n21874), .ip2(n21868), .op(n21869) );
  xor2_1 U24604 ( .ip1(n21870), .ip2(n21869), .op(n21871) );
  nand2_1 U24605 ( .ip1(n21944), .ip2(n21871), .op(n21872) );
  nand2_1 U24606 ( .ip1(n21873), .ip2(n21872), .op(n8550) );
  nand2_1 U24607 ( .ip1(\pipeline/md/a [53]), .ip2(n21884), .op(n21883) );
  inv_1 U24608 ( .ip(n21874), .op(n21876) );
  nor2_1 U24609 ( .ip1(n21876), .ip2(n21875), .op(n21880) );
  nand2_1 U24610 ( .ip1(n21878), .ip2(n21877), .op(n21879) );
  xor2_1 U24611 ( .ip1(n21880), .ip2(n21879), .op(n21881) );
  nand2_1 U24612 ( .ip1(n21944), .ip2(n21881), .op(n21882) );
  nand2_1 U24613 ( .ip1(n21883), .ip2(n21882), .op(n8549) );
  nand2_1 U24614 ( .ip1(\pipeline/md/a [54]), .ip2(n21884), .op(n21890) );
  nand2_1 U24615 ( .ip1(n21891), .ip2(n21885), .op(n21886) );
  xor2_1 U24616 ( .ip1(n21887), .ip2(n21886), .op(n21888) );
  nand2_1 U24617 ( .ip1(n21944), .ip2(n21888), .op(n21889) );
  nand2_1 U24618 ( .ip1(n21890), .ip2(n21889), .op(n8548) );
  nand2_1 U24619 ( .ip1(\pipeline/md/a [55]), .ip2(n21947), .op(n21901) );
  inv_1 U24620 ( .ip(n21891), .op(n21893) );
  nor2_1 U24621 ( .ip1(n21893), .ip2(n21892), .op(n21898) );
  inv_1 U24622 ( .ip(n21894), .op(n21895) );
  nand2_1 U24623 ( .ip1(n21896), .ip2(n21895), .op(n21897) );
  xor2_1 U24624 ( .ip1(n21898), .ip2(n21897), .op(n21899) );
  nand2_1 U24625 ( .ip1(n21944), .ip2(n21899), .op(n21900) );
  nand2_1 U24626 ( .ip1(n21901), .ip2(n21900), .op(n8547) );
  xor2_1 U24627 ( .ip1(\pipeline/md/b [56]), .ip2(n21909), .op(n21902) );
  nor2_1 U24628 ( .ip1(\pipeline/md/a [56]), .ip2(n21902), .op(n21903) );
  nand2_1 U24629 ( .ip1(n21944), .ip2(n21903), .op(n21914) );
  inv_1 U24630 ( .ip(n21904), .op(n21908) );
  nor2_1 U24631 ( .ip1(n21905), .ip2(n21910), .op(n21906) );
  nor2_1 U24632 ( .ip1(n21909), .ip2(n21906), .op(n21907) );
  not_ab_or_c_or_d U24633 ( .ip1(n21909), .ip2(n21908), .ip3(n21907), .ip4(
        n22665), .op(n21912) );
  nor2_1 U24634 ( .ip1(n21910), .ip2(n14770), .op(n21911) );
  nor2_1 U24635 ( .ip1(n21912), .ip2(n21911), .op(n21913) );
  nand2_1 U24636 ( .ip1(n21914), .ip2(n21913), .op(n8546) );
  xor2_1 U24637 ( .ip1(\pipeline/md/b [57]), .ip2(n21917), .op(n21915) );
  nor2_1 U24638 ( .ip1(\pipeline/md/a [57]), .ip2(n21915), .op(n21916) );
  nand2_1 U24639 ( .ip1(n21944), .ip2(n21916), .op(n21926) );
  inv_1 U24640 ( .ip(n21917), .op(n21921) );
  nand2_1 U24641 ( .ip1(\pipeline/md/b [57]), .ip2(\pipeline/md/a [57]), .op(
        n21920) );
  nor2_1 U24642 ( .ip1(n21918), .ip2(n21921), .op(n21919) );
  not_ab_or_c_or_d U24643 ( .ip1(n21921), .ip2(n21920), .ip3(n21919), .ip4(
        n22665), .op(n21924) );
  nor2_1 U24644 ( .ip1(n21922), .ip2(n14770), .op(n21923) );
  nor2_1 U24645 ( .ip1(n21924), .ip2(n21923), .op(n21925) );
  nand2_1 U24646 ( .ip1(n21926), .ip2(n21925), .op(n8545) );
  xor2_1 U24647 ( .ip1(\pipeline/md/b [58]), .ip2(n21937), .op(n21927) );
  nand2_1 U24648 ( .ip1(n20310), .ip2(n21927), .op(n21928) );
  nand2_1 U24649 ( .ip1(n14770), .ip2(n21928), .op(n21929) );
  nand2_1 U24650 ( .ip1(\pipeline/md/a [58]), .ip2(n21929), .op(n21933) );
  nor2_1 U24651 ( .ip1(\pipeline/md/b [58]), .ip2(\pipeline/md/a [58]), .op(
        n21930) );
  mux2_1 U24652 ( .ip1(n21930), .ip2(n21940), .s(n21937), .op(n21931) );
  nand2_1 U24653 ( .ip1(n21944), .ip2(n21931), .op(n21932) );
  nand2_1 U24654 ( .ip1(n21933), .ip2(n21932), .op(n8544) );
  nand2_1 U24655 ( .ip1(\pipeline/md/a [59]), .ip2(n21947), .op(n21946) );
  nor2_1 U24656 ( .ip1(n21935), .ip2(n21934), .op(n21942) );
  inv_1 U24657 ( .ip(n21936), .op(n21938) );
  nor2_1 U24658 ( .ip1(n21938), .ip2(n21937), .op(n21939) );
  nor2_1 U24659 ( .ip1(n21940), .ip2(n21939), .op(n21941) );
  xor2_1 U24660 ( .ip1(n21942), .ip2(n21941), .op(n21943) );
  nand2_1 U24661 ( .ip1(n21944), .ip2(n21943), .op(n21945) );
  nand2_1 U24662 ( .ip1(n21946), .ip2(n21945), .op(n8543) );
  nand2_1 U24663 ( .ip1(n21947), .ip2(\pipeline/md/a [62]), .op(n21954) );
  fulladder U24664 ( .a(n21949), .b(\pipeline/md/b [61]), .ci(n21948), .co(
        n21950), .s(n21736) );
  fulladder U24665 ( .a(\pipeline/md/b [62]), .b(n21951), .ci(n21950), .co(), 
        .s(n21952) );
  or2_1 U24666 ( .ip1(n21952), .ip2(n21730), .op(n21953) );
  nand2_1 U24667 ( .ip1(n21954), .ip2(n21953), .op(n8540) );
  nor4_1 U24668 ( .ip1(\pipeline/md_resp_result [24]), .ip2(n21979), .ip3(
        n15245), .ip4(n22755), .op(n21976) );
  nand2_1 U24669 ( .ip1(\pipeline/md/negate_output ), .ip2(n21955), .op(n21956) );
  nor2_1 U24670 ( .ip1(n21959), .ip2(n21956), .op(n21964) );
  nor2_1 U24671 ( .ip1(n21958), .ip2(n21957), .op(n21962) );
  nor2_1 U24672 ( .ip1(n21960), .ip2(n21959), .op(n21961) );
  nor2_1 U24673 ( .ip1(n21962), .ip2(n21961), .op(n21963) );
  nor2_1 U24674 ( .ip1(n21964), .ip2(n21963), .op(n21974) );
  inv_1 U24675 ( .ip(n21969), .op(n21965) );
  nor3_1 U24676 ( .ip1(\pipeline/md/result [56]), .ip2(n21966), .ip3(n21965), 
        .op(n21971) );
  inv_1 U24677 ( .ip(\pipeline/md/result [56]), .op(n21968) );
  not_ab_or_c_or_d U24678 ( .ip1(\pipeline/md/negate_output ), .ip2(n21969), 
        .ip3(n21968), .ip4(n21967), .op(n21970) );
  nor3_1 U24679 ( .ip1(n21972), .ip2(n21971), .ip3(n21970), .op(n21973) );
  nor2_1 U24680 ( .ip1(n21974), .ip2(n21973), .op(n21975) );
  not_ab_or_c_or_d U24681 ( .ip1(n21978), .ip2(n21977), .ip3(n21976), .ip4(
        n21975), .op(n21984) );
  or2_1 U24682 ( .ip1(n21979), .ip2(n15245), .op(n21980) );
  nand2_1 U24683 ( .ip1(n14765), .ip2(n21980), .op(n21981) );
  nand2_1 U24684 ( .ip1(n22738), .ip2(n21981), .op(n21982) );
  nand2_1 U24685 ( .ip1(\pipeline/md_resp_result [24]), .ip2(n21982), .op(
        n21983) );
  nand2_1 U24686 ( .ip1(n21984), .ip2(n21983), .op(n8610) );
  mux2_1 U24687 ( .ip1(\pipeline/csr_rdata_WB [24]), .ip2(n21985), .s(n17429), 
        .op(n8782) );
  nand2_1 U24688 ( .ip1(\pipeline/PC_IF [31]), .ip2(n21996), .op(n21986) );
  nand2_1 U24689 ( .ip1(n21987), .ip2(n21986), .op(n8428) );
  nand2_1 U24690 ( .ip1(\pipeline/PC_IF [31]), .ip2(n21988), .op(n21990) );
  nand2_1 U24691 ( .ip1(\pipeline/PC_DX [31]), .ip2(n21999), .op(n21989) );
  nand2_1 U24692 ( .ip1(n21990), .ip2(n21989), .op(n8427) );
  nor2_1 U24693 ( .ip1(n21992), .ip2(n21991), .op(n21993) );
  nor2_1 U24694 ( .ip1(n21994), .ip2(n21993), .op(imem_haddr[1]) );
  nand2_1 U24695 ( .ip1(n21995), .ip2(imem_haddr[1]), .op(n21998) );
  nand2_1 U24696 ( .ip1(\pipeline/PC_IF [1]), .ip2(n21996), .op(n21997) );
  nand2_1 U24697 ( .ip1(n21998), .ip2(n21997), .op(n8488) );
  nand2_1 U24698 ( .ip1(\pipeline/PC_IF [1]), .ip2(n22048), .op(n22001) );
  nand2_1 U24699 ( .ip1(\pipeline/PC_DX [1]), .ip2(n21999), .op(n22000) );
  nand2_1 U24700 ( .ip1(n22001), .ip2(n22000), .op(n8487) );
  mux2_1 U24701 ( .ip1(\pipeline/PC_WB [1]), .ip2(\pipeline/PC_DX [1]), .s(
        n20389), .op(n8902) );
  xor2_1 U24702 ( .ip1(\pipeline/csr/time_full [0]), .ip2(
        \pipeline/csr/time_full [1]), .op(n22004) );
  inv_1 U24703 ( .ip(n22002), .op(n22003) );
  nand2_1 U24704 ( .ip1(n22004), .ip2(n22003), .op(n22007) );
  nand2_1 U24705 ( .ip1(n22005), .ip2(n22129), .op(n22006) );
  nand2_1 U24706 ( .ip1(n22007), .ip2(n22006), .op(\pipeline/csr/N1938 ) );
  nand2_1 U24707 ( .ip1(n22008), .ip2(n22129), .op(n22012) );
  xor2_1 U24708 ( .ip1(\pipeline/csr/mtime_full [0]), .ip2(
        \pipeline/csr/mtime_full [1]), .op(n22010) );
  nand2_1 U24709 ( .ip1(n22010), .ip2(n22009), .op(n22011) );
  nand2_1 U24710 ( .ip1(n22012), .ip2(n22011), .op(\pipeline/csr/N2082 ) );
  nand2_1 U24711 ( .ip1(n22013), .ip2(\pipeline/csr/mscratch [1]), .op(n22016)
         );
  nand2_1 U24712 ( .ip1(n22014), .ip2(n22129), .op(n22015) );
  nand2_1 U24713 ( .ip1(n22016), .ip2(n22015), .op(n9927) );
  nand2_1 U24714 ( .ip1(n22372), .ip2(\pipeline/csr/from_host [1]), .op(n22018) );
  nand2_1 U24715 ( .ip1(n22373), .ip2(n22129), .op(n22017) );
  nand2_1 U24716 ( .ip1(n22018), .ip2(n22017), .op(n9959) );
  nand2_1 U24717 ( .ip1(n22378), .ip2(n22129), .op(n22020) );
  nand2_1 U24718 ( .ip1(n22376), .ip2(\pipeline/csr/to_host [1]), .op(n22019)
         );
  nand2_1 U24719 ( .ip1(n22020), .ip2(n22019), .op(n8771) );
  nand2_1 U24720 ( .ip1(n22021), .ip2(n22129), .op(n22025) );
  xor2_1 U24721 ( .ip1(\pipeline/csr/cycle_full [0]), .ip2(
        \pipeline/csr/cycle_full [1]), .op(n22023) );
  nand2_1 U24722 ( .ip1(n22023), .ip2(n22022), .op(n22024) );
  nand2_1 U24723 ( .ip1(n22025), .ip2(n22024), .op(\pipeline/csr/N1874 ) );
  nand2_1 U24724 ( .ip1(n22363), .ip2(\pipeline/csr/mtimecmp [1]), .op(n22027)
         );
  nand2_1 U24725 ( .ip1(n22365), .ip2(n22129), .op(n22026) );
  nand2_1 U24726 ( .ip1(n22027), .ip2(n22026), .op(n10021) );
  nand2_1 U24727 ( .ip1(n22356), .ip2(\pipeline/csr/mie [1]), .op(n22029) );
  nand2_1 U24728 ( .ip1(n22357), .ip2(n22129), .op(n22028) );
  nand2_1 U24729 ( .ip1(n22029), .ip2(n22028), .op(n10059) );
  nor2_1 U24730 ( .ip1(n22261), .ip2(n22305), .op(n22032) );
  not_ab_or_c_or_d U24731 ( .ip1(n22291), .ip2(n22030), .ip3(n22294), .ip4(
        n22308), .op(n22031) );
  or2_1 U24732 ( .ip1(n22032), .ip2(n22031), .op(\pipeline/csr/N1906 ) );
  nor2_1 U24733 ( .ip1(n22033), .ip2(n22036), .op(n22035) );
  not_ab_or_c_or_d U24734 ( .ip1(\pipeline/csr/priv_stack [4]), .ip2(n22036), 
        .ip3(n22035), .ip4(n22034), .op(n22039) );
  nor2_1 U24735 ( .ip1(\pipeline/prv [0]), .ip2(n22037), .op(n22038) );
  nor2_1 U24736 ( .ip1(n22039), .ip2(n22038), .op(n10026) );
  nand2_1 U24737 ( .ip1(n22048), .ip2(imem_rdata[25]), .op(n22041) );
  nand2_1 U24738 ( .ip1(\pipeline/inst_DX [25]), .ip2(n22049), .op(n22040) );
  nand2_1 U24739 ( .ip1(n22041), .ip2(n22040), .op(n8510) );
  nand2_1 U24740 ( .ip1(n22042), .ip2(n17429), .op(n22045) );
  nand2_1 U24741 ( .ip1(\pipeline/ctrl/uses_md_WB ), .ip2(n22043), .op(n22044)
         );
  nand2_1 U24742 ( .ip1(n22045), .ip2(n22044), .op(n8493) );
  inv_1 U24743 ( .ip(n22046), .op(n22047) );
  nor2_1 U24744 ( .ip1(n22047), .ip2(n21582), .op(n8499) );
  nand2_1 U24745 ( .ip1(n22048), .ip2(imem_rdata[30]), .op(n22051) );
  nand2_1 U24746 ( .ip1(\pipeline/inst_DX [30]), .ip2(n22049), .op(n22050) );
  nand2_1 U24747 ( .ip1(n22051), .ip2(n22050), .op(n8505) );
  mux2_1 U24748 ( .ip1(\pipeline/store_data_WB [24]), .ip2(n21278), .s(n19498), 
        .op(n8815) );
  mux2_1 U24749 ( .ip1(\pipeline/store_data_WB [25]), .ip2(n21282), .s(n19498), 
        .op(n8814) );
  mux2_1 U24750 ( .ip1(dmem_hwdata[2]), .ip2(n22057), .s(n20389), .op(n8837)
         );
  mux2_1 U24751 ( .ip1(\pipeline/store_data_WB [26]), .ip2(n21281), .s(n17777), 
        .op(n8813) );
  mux2_1 U24752 ( .ip1(\pipeline/store_data_WB [27]), .ip2(n21277), .s(n17429), 
        .op(n8812) );
  mux2_1 U24753 ( .ip1(\pipeline/store_data_WB [28]), .ip2(n21276), .s(n22067), 
        .op(n8811) );
  inv_1 U24754 ( .ip(\pipeline/dmem_type_WB [2]), .op(n22070) );
  nand2_1 U24755 ( .ip1(n22071), .ip2(n22070), .op(n22079) );
  nand2_1 U24756 ( .ip1(\pipeline/store_data_WB [8]), .ip2(n22079), .op(n22072) );
  inv_1 U24757 ( .ip(n22079), .op(n22080) );
  nand2_1 U24758 ( .ip1(dmem_hwdata[0]), .ip2(n22080), .op(n22322) );
  nand2_1 U24759 ( .ip1(n22072), .ip2(n22322), .op(dmem_hwdata[8]) );
  nand2_1 U24760 ( .ip1(\pipeline/store_data_WB [9]), .ip2(n22079), .op(n22073) );
  nand2_1 U24761 ( .ip1(dmem_hwdata[1]), .ip2(n22080), .op(n22326) );
  nand2_1 U24762 ( .ip1(n22073), .ip2(n22326), .op(dmem_hwdata[9]) );
  nand2_1 U24763 ( .ip1(\pipeline/store_data_WB [10]), .ip2(n22079), .op(
        n22074) );
  nand2_1 U24764 ( .ip1(dmem_hwdata[2]), .ip2(n22080), .op(n22329) );
  nand2_1 U24765 ( .ip1(n22074), .ip2(n22329), .op(dmem_hwdata[10]) );
  nand2_1 U24766 ( .ip1(\pipeline/store_data_WB [11]), .ip2(n22079), .op(
        n22075) );
  nand2_1 U24767 ( .ip1(dmem_hwdata[3]), .ip2(n22080), .op(n22332) );
  nand2_1 U24768 ( .ip1(n22075), .ip2(n22332), .op(dmem_hwdata[11]) );
  nand2_1 U24769 ( .ip1(\pipeline/store_data_WB [12]), .ip2(n22079), .op(
        n22076) );
  nand2_1 U24770 ( .ip1(dmem_hwdata[4]), .ip2(n22080), .op(n22335) );
  nand2_1 U24771 ( .ip1(n22076), .ip2(n22335), .op(dmem_hwdata[12]) );
  nand2_1 U24772 ( .ip1(\pipeline/store_data_WB [13]), .ip2(n22079), .op(
        n22077) );
  nand2_1 U24773 ( .ip1(dmem_hwdata[5]), .ip2(n22080), .op(n22338) );
  nand2_1 U24774 ( .ip1(n22077), .ip2(n22338), .op(dmem_hwdata[13]) );
  nand2_1 U24775 ( .ip1(\pipeline/store_data_WB [14]), .ip2(n22079), .op(
        n22078) );
  nand2_1 U24776 ( .ip1(dmem_hwdata[6]), .ip2(n22080), .op(n22341) );
  nand2_1 U24777 ( .ip1(n22078), .ip2(n22341), .op(dmem_hwdata[14]) );
  nand2_1 U24778 ( .ip1(\pipeline/store_data_WB [15]), .ip2(n22079), .op(
        n22081) );
  nand2_1 U24779 ( .ip1(dmem_hwdata[7]), .ip2(n22080), .op(n22346) );
  nand2_1 U24780 ( .ip1(n22081), .ip2(n22346), .op(dmem_hwdata[15]) );
  mux2_1 U24781 ( .ip1(\pipeline/store_data_WB [16]), .ip2(dmem_hwdata[0]), 
        .s(n22087), .op(dmem_hwdata[16]) );
  mux2_1 U24782 ( .ip1(\pipeline/store_data_WB [17]), .ip2(n17387), .s(n17429), 
        .op(n8822) );
  mux2_1 U24783 ( .ip1(\pipeline/store_data_WB [17]), .ip2(dmem_hwdata[1]), 
        .s(n22087), .op(dmem_hwdata[17]) );
  mux2_1 U24784 ( .ip1(\pipeline/store_data_WB [18]), .ip2(dmem_hwdata[2]), 
        .s(n22087), .op(dmem_hwdata[18]) );
  mux2_1 U24785 ( .ip1(\pipeline/store_data_WB [19]), .ip2(dmem_hwdata[3]), 
        .s(n22087), .op(dmem_hwdata[19]) );
  mux2_1 U24786 ( .ip1(\pipeline/store_data_WB [20]), .ip2(dmem_hwdata[4]), 
        .s(n22087), .op(dmem_hwdata[20]) );
  mux2_1 U24787 ( .ip1(\pipeline/store_data_WB [21]), .ip2(dmem_hwdata[5]), 
        .s(n22087), .op(dmem_hwdata[21]) );
  mux2_1 U24788 ( .ip1(\pipeline/store_data_WB [22]), .ip2(n22086), .s(n17429), 
        .op(n8817) );
  mux2_1 U24789 ( .ip1(\pipeline/store_data_WB [22]), .ip2(dmem_hwdata[6]), 
        .s(n22087), .op(dmem_hwdata[22]) );
  mux2_1 U24790 ( .ip1(\pipeline/store_data_WB [23]), .ip2(dmem_hwdata[7]), 
        .s(n22087), .op(dmem_hwdata[23]) );
  nand2_1 U24791 ( .ip1(\pipeline/csr/mie [5]), .ip2(n22356), .op(n22089) );
  nand2_1 U24792 ( .ip1(n22357), .ip2(n22145), .op(n22088) );
  nand2_1 U24793 ( .ip1(n22089), .ip2(n22088), .op(n10055) );
  and2_1 U24794 ( .ip1(n22091), .ip2(n22090), .op(n22866) );
  or2_1 U24795 ( .ip1(n22092), .ip2(n22098), .op(n22118) );
  inv_1 U24796 ( .ip(n22118), .op(n22107) );
  nor2_1 U24797 ( .ip1(n22107), .ip2(n22093), .op(n22117) );
  nor4_1 U24798 ( .ip1(\pipeline/inst_DX [23]), .ip2(\pipeline/inst_DX [22]), 
        .ip3(n22094), .ip4(n22100), .op(n22095) );
  not_ab_or_c_or_d U24799 ( .ip1(n22098), .ip2(n22097), .ip3(n22096), .ip4(
        n22095), .op(n22115) );
  inv_1 U24800 ( .ip(n22099), .op(n22102) );
  inv_1 U24801 ( .ip(n22100), .op(n22101) );
  not_ab_or_c_or_d U24802 ( .ip1(n22104), .ip2(n22103), .ip3(n22102), .ip4(
        n22101), .op(n22106) );
  nand3_1 U24803 ( .ip1(n22107), .ip2(n22106), .ip3(n22105), .op(n22108) );
  nand2_1 U24804 ( .ip1(n22109), .ip2(n22108), .op(n22114) );
  inv_1 U24805 ( .ip(n22110), .op(n22111) );
  nand2_1 U24806 ( .ip1(n22112), .ip2(n22111), .op(n22113) );
  nand3_1 U24807 ( .ip1(n22115), .ip2(n22114), .ip3(n22113), .op(n22116) );
  not_ab_or_c_or_d U24808 ( .ip1(n22119), .ip2(n22118), .ip3(n22117), .ip4(
        n22116), .op(n10142) );
  nor2_1 U24809 ( .ip1(\pipeline/prv [1]), .ip2(n22121), .op(n22123) );
  not_ab_or_c_or_d U24810 ( .ip1(\pipeline/prv [1]), .ip2(n22121), .ip3(
        \pipeline/prv [0]), .ip4(n22120), .op(n22122) );
  or2_1 U24811 ( .ip1(n22123), .ip2(n22122), .op(n10143) );
  not_ab_or_c_or_d U24814 ( .ip1(n22125), .ip2(n22124), .ip3(n22247), .ip4(
        n22130), .op(n22128) );
  inv_1 U24815 ( .ip(n22377), .op(n22126) );
  nor2_1 U24816 ( .ip1(n22126), .ip2(n22244), .op(n22127) );
  or2_1 U24817 ( .ip1(n22128), .ip2(n22127), .op(\pipeline/csr/N2113 ) );
  nand2_1 U24818 ( .ip1(n22235), .ip2(n22129), .op(n22133) );
  or2_1 U24819 ( .ip1(\pipeline/csr/mtime_full [33]), .ip2(n22130), .op(n22131) );
  nand3_1 U24820 ( .ip1(n22136), .ip2(n22131), .ip3(n18449), .op(n22132) );
  nand2_1 U24821 ( .ip1(n22133), .ip2(n22132), .op(\pipeline/csr/N2114 ) );
  nor2_1 U24822 ( .ip1(n22134), .ip2(n22244), .op(n22139) );
  not_ab_or_c_or_d U24823 ( .ip1(n22137), .ip2(n22136), .ip3(n22247), .ip4(
        n22135), .op(n22138) );
  or2_1 U24824 ( .ip1(n22139), .ip2(n22138), .op(\pipeline/csr/N2115 ) );
  inv_1 U24825 ( .ip(n22360), .op(n22140) );
  nor2_1 U24826 ( .ip1(n22140), .ip2(n22244), .op(n22144) );
  not_ab_or_c_or_d U24827 ( .ip1(n22142), .ip2(n22141), .ip3(n22247), .ip4(
        n22146), .op(n22143) );
  or2_1 U24828 ( .ip1(n22144), .ip2(n22143), .op(\pipeline/csr/N2117 ) );
  nand2_1 U24829 ( .ip1(n22235), .ip2(n22145), .op(n22149) );
  or2_1 U24830 ( .ip1(\pipeline/csr/mtime_full [37]), .ip2(n22146), .op(n22147) );
  nand3_1 U24831 ( .ip1(n22152), .ip2(n22147), .ip3(n18449), .op(n22148) );
  nand2_1 U24832 ( .ip1(n22149), .ip2(n22148), .op(\pipeline/csr/N2118 ) );
  inv_1 U24833 ( .ip(n22364), .op(n22150) );
  nor2_1 U24834 ( .ip1(n22150), .ip2(n22244), .op(n22155) );
  not_ab_or_c_or_d U24835 ( .ip1(n22153), .ip2(n22152), .ip3(n22247), .ip4(
        n22151), .op(n22154) );
  or2_1 U24836 ( .ip1(n22155), .ip2(n22154), .op(\pipeline/csr/N2119 ) );
  nand2_1 U24837 ( .ip1(n22235), .ip2(n22156), .op(n22160) );
  or2_1 U24838 ( .ip1(\pipeline/csr/mtime_full [43]), .ip2(n22157), .op(n22158) );
  nand3_1 U24839 ( .ip1(n22162), .ip2(n22158), .ip3(n18449), .op(n22159) );
  nand2_1 U24840 ( .ip1(n22160), .ip2(n22159), .op(\pipeline/csr/N2124 ) );
  nor2_1 U24841 ( .ip1(n22161), .ip2(n22244), .op(n22165) );
  not_ab_or_c_or_d U24842 ( .ip1(n22163), .ip2(n22162), .ip3(n22247), .ip4(
        n22167), .op(n22164) );
  or2_1 U24843 ( .ip1(n22165), .ip2(n22164), .op(\pipeline/csr/N2125 ) );
  nand2_1 U24844 ( .ip1(n22235), .ip2(n22166), .op(n22170) );
  or2_1 U24845 ( .ip1(\pipeline/csr/mtime_full [45]), .ip2(n22167), .op(n22168) );
  nand3_1 U24846 ( .ip1(n22173), .ip2(n22168), .ip3(n18449), .op(n22169) );
  nand2_1 U24847 ( .ip1(n22170), .ip2(n22169), .op(\pipeline/csr/N2126 ) );
  inv_1 U24848 ( .ip(n22171), .op(n22172) );
  nor2_1 U24849 ( .ip1(n22172), .ip2(n22244), .op(n22176) );
  not_ab_or_c_or_d U24850 ( .ip1(n22174), .ip2(n22173), .ip3(n22247), .ip4(
        n22178), .op(n22175) );
  or2_1 U24851 ( .ip1(n22176), .ip2(n22175), .op(\pipeline/csr/N2127 ) );
  nand2_1 U24852 ( .ip1(n22235), .ip2(n22177), .op(n22182) );
  or2_1 U24853 ( .ip1(\pipeline/csr/mtime_full [47]), .ip2(n22178), .op(n22179) );
  nand3_1 U24854 ( .ip1(n22180), .ip2(n22179), .ip3(n18449), .op(n22181) );
  nand2_1 U24855 ( .ip1(n22182), .ip2(n22181), .op(\pipeline/csr/N2128 ) );
  nand2_1 U24856 ( .ip1(n22235), .ip2(n22183), .op(n22188) );
  or2_1 U24857 ( .ip1(\pipeline/csr/mtime_full [49]), .ip2(n22184), .op(n22185) );
  nand3_1 U24858 ( .ip1(n22186), .ip2(n22185), .ip3(n18449), .op(n22187) );
  nand2_1 U24859 ( .ip1(n22188), .ip2(n22187), .op(\pipeline/csr/N2130 ) );
  nand2_1 U24860 ( .ip1(n22235), .ip2(n22189), .op(n22193) );
  or2_1 U24861 ( .ip1(\pipeline/csr/mtime_full [51]), .ip2(n22190), .op(n22191) );
  nand3_1 U24862 ( .ip1(n22195), .ip2(n22191), .ip3(n18449), .op(n22192) );
  nand2_1 U24863 ( .ip1(n22193), .ip2(n22192), .op(\pipeline/csr/N2132 ) );
  nor2_1 U24864 ( .ip1(n22194), .ip2(n22244), .op(n22198) );
  not_ab_or_c_or_d U24865 ( .ip1(n22196), .ip2(n22195), .ip3(n22247), .ip4(
        n22199), .op(n22197) );
  or2_1 U24866 ( .ip1(n22198), .ip2(n22197), .op(\pipeline/csr/N2133 ) );
  nand2_1 U24867 ( .ip1(n22235), .ip2(n22368), .op(n22202) );
  or2_1 U24868 ( .ip1(\pipeline/csr/mtime_full [53]), .ip2(n22199), .op(n22200) );
  nand3_1 U24869 ( .ip1(n22204), .ip2(n22200), .ip3(n18449), .op(n22201) );
  nand2_1 U24870 ( .ip1(n22202), .ip2(n22201), .op(\pipeline/csr/N2134 ) );
  nor2_1 U24871 ( .ip1(n22203), .ip2(n22244), .op(n22207) );
  not_ab_or_c_or_d U24872 ( .ip1(n22205), .ip2(n22204), .ip3(n22247), .ip4(
        n22208), .op(n22206) );
  or2_1 U24873 ( .ip1(n22207), .ip2(n22206), .op(\pipeline/csr/N2135 ) );
  nand2_1 U24874 ( .ip1(n22235), .ip2(n22274), .op(n22211) );
  or2_1 U24875 ( .ip1(\pipeline/csr/mtime_full [55]), .ip2(n22208), .op(n22209) );
  nand3_1 U24876 ( .ip1(n22213), .ip2(n22209), .ip3(n18449), .op(n22210) );
  nand2_1 U24877 ( .ip1(n22211), .ip2(n22210), .op(\pipeline/csr/N2136 ) );
  nor2_1 U24878 ( .ip1(n22212), .ip2(n22244), .op(n22216) );
  not_ab_or_c_or_d U24879 ( .ip1(n22214), .ip2(n22213), .ip3(n22247), .ip4(
        n22218), .op(n22215) );
  or2_1 U24880 ( .ip1(n22216), .ip2(n22215), .op(\pipeline/csr/N2137 ) );
  nand2_1 U24881 ( .ip1(n22235), .ip2(n22217), .op(n22221) );
  or2_1 U24882 ( .ip1(\pipeline/csr/mtime_full [57]), .ip2(n22218), .op(n22219) );
  nand3_1 U24883 ( .ip1(n22225), .ip2(n22219), .ip3(n18449), .op(n22220) );
  nand2_1 U24884 ( .ip1(n22221), .ip2(n22220), .op(\pipeline/csr/N2138 ) );
  inv_1 U24885 ( .ip(n22222), .op(n22223) );
  nor2_1 U24886 ( .ip1(n22223), .ip2(n22244), .op(n22228) );
  not_ab_or_c_or_d U24887 ( .ip1(n22226), .ip2(n22225), .ip3(n22247), .ip4(
        n22224), .op(n22227) );
  or2_1 U24888 ( .ip1(n22228), .ip2(n22227), .op(\pipeline/csr/N2139 ) );
  nor2_1 U24889 ( .ip1(n22229), .ip2(n22244), .op(n22233) );
  nor2_1 U24890 ( .ip1(n22231), .ip2(n22230), .op(n22236) );
  not_ab_or_c_or_d U24891 ( .ip1(n22231), .ip2(n22230), .ip3(n22247), .ip4(
        n22236), .op(n22232) );
  or2_1 U24892 ( .ip1(n22233), .ip2(n22232), .op(\pipeline/csr/N2141 ) );
  nand2_1 U24893 ( .ip1(n22235), .ip2(n22234), .op(n22239) );
  nand2_1 U24894 ( .ip1(\pipeline/csr/mtime_full [61]), .ip2(n22236), .op(
        n22240) );
  or2_1 U24895 ( .ip1(\pipeline/csr/mtime_full [61]), .ip2(n22236), .op(n22237) );
  nand3_1 U24896 ( .ip1(n22240), .ip2(n22237), .ip3(n18449), .op(n22238) );
  nand2_1 U24897 ( .ip1(n22239), .ip2(n22238), .op(\pipeline/csr/N2142 ) );
  nor2_1 U24898 ( .ip1(n22258), .ip2(n22244), .op(n22243) );
  inv_1 U24899 ( .ip(\pipeline/csr/mtime_full [62]), .op(n22241) );
  nor2_1 U24900 ( .ip1(n22241), .ip2(n22240), .op(n22248) );
  not_ab_or_c_or_d U24901 ( .ip1(n22241), .ip2(n22240), .ip3(n22247), .ip4(
        n22248), .op(n22242) );
  or2_1 U24902 ( .ip1(n22243), .ip2(n22242), .op(\pipeline/csr/N2143 ) );
  nor2_1 U24903 ( .ip1(n22245), .ip2(n22244), .op(n22250) );
  nor2_1 U24904 ( .ip1(\pipeline/csr/mtime_full [63]), .ip2(n22248), .op(
        n22246) );
  not_ab_or_c_or_d U24905 ( .ip1(\pipeline/csr/mtime_full [63]), .ip2(n22248), 
        .ip3(n22247), .ip4(n22246), .op(n22249) );
  or2_1 U24906 ( .ip1(n22250), .ip2(n22249), .op(\pipeline/csr/N2144 ) );
  xor2_1 U24907 ( .ip1(\pipeline/csr/time_full [30]), .ip2(n22251), .op(n22253) );
  nand2_1 U24908 ( .ip1(n22253), .ip2(n22252), .op(n22260) );
  nor2_1 U24909 ( .ip1(n22254), .ip2(n22253), .op(n22256) );
  ab_or_c_or_d U24910 ( .ip1(n22258), .ip2(n22257), .ip3(n22256), .ip4(n22255), 
        .op(n22259) );
  nand2_1 U24911 ( .ip1(n22260), .ip2(n22259), .op(\pipeline/csr/N1967 ) );
  nor2_1 U24912 ( .ip1(n22261), .ip2(n22267), .op(n22266) );
  not_ab_or_c_or_d U24913 ( .ip1(n22264), .ip2(n22263), .ip3(n22276), .ip4(
        n22262), .op(n22265) );
  or2_1 U24914 ( .ip1(n22266), .ip2(n22265), .op(\pipeline/csr/N1970 ) );
  nor2_1 U24915 ( .ip1(n22268), .ip2(n22267), .op(n22273) );
  not_ab_or_c_or_d U24916 ( .ip1(n22271), .ip2(n22270), .ip3(n22276), .ip4(
        n22269), .op(n22272) );
  or2_1 U24917 ( .ip1(n22273), .ip2(n22272), .op(\pipeline/csr/N1972 ) );
  nand2_1 U24918 ( .ip1(n22282), .ip2(n22274), .op(n22280) );
  ab_or_c_or_d U24919 ( .ip1(n22278), .ip2(n22277), .ip3(n22276), .ip4(n22275), 
        .op(n22279) );
  nand2_1 U24920 ( .ip1(n22280), .ip2(n22279), .op(\pipeline/csr/N1992 ) );
  nand2_1 U24921 ( .ip1(n22282), .ip2(n22281), .op(n22288) );
  or2_1 U24922 ( .ip1(\pipeline/csr/time_full [60]), .ip2(n22283), .op(n22285)
         );
  nand3_1 U24923 ( .ip1(n22286), .ip2(n22285), .ip3(n22284), .op(n22287) );
  nand2_1 U24924 ( .ip1(n22288), .ip2(n22287), .op(\pipeline/csr/N1997 ) );
  or2_1 U24925 ( .ip1(\pipeline/csr/cycle_full [32]), .ip2(n22289), .op(n22290) );
  nand3_1 U24926 ( .ip1(n22291), .ip2(n22290), .ip3(n22316), .op(n22293) );
  nand2_1 U24927 ( .ip1(n22314), .ip2(n22377), .op(n22292) );
  nand2_1 U24928 ( .ip1(n22293), .ip2(n22292), .op(\pipeline/csr/N1905 ) );
  nand2_1 U24929 ( .ip1(n22314), .ip2(n22351), .op(n22298) );
  or2_1 U24930 ( .ip1(\pipeline/csr/cycle_full [34]), .ip2(n22294), .op(n22295) );
  nand3_1 U24931 ( .ip1(n22296), .ip2(n22295), .ip3(n22316), .op(n22297) );
  nand2_1 U24932 ( .ip1(n22298), .ip2(n22297), .op(\pipeline/csr/N1907 ) );
  nor2_1 U24933 ( .ip1(n22299), .ip2(n22305), .op(n22304) );
  not_ab_or_c_or_d U24934 ( .ip1(n22302), .ip2(n22301), .ip3(n22308), .ip4(
        n22300), .op(n22303) );
  or2_1 U24935 ( .ip1(n22304), .ip2(n22303), .op(\pipeline/csr/N1928 ) );
  nor2_1 U24936 ( .ip1(n22306), .ip2(n22305), .op(n22312) );
  not_ab_or_c_or_d U24937 ( .ip1(n22310), .ip2(n22309), .ip3(n22308), .ip4(
        n22307), .op(n22311) );
  or2_1 U24938 ( .ip1(n22312), .ip2(n22311), .op(\pipeline/csr/N1930 ) );
  nand2_1 U24939 ( .ip1(n22314), .ip2(n22313), .op(n22320) );
  or2_1 U24940 ( .ip1(\pipeline/csr/cycle_full [62]), .ip2(n22315), .op(n22317) );
  nand3_1 U24941 ( .ip1(n22318), .ip2(n22317), .ip3(n22316), .op(n22319) );
  nand2_1 U24942 ( .ip1(n22320), .ip2(n22319), .op(\pipeline/csr/N1935 ) );
  inv_1 U24943 ( .ip(n22321), .op(n22343) );
  nand2_1 U24944 ( .ip1(n22343), .ip2(\pipeline/store_data_WB [8]), .op(n22324) );
  nand2_1 U24945 ( .ip1(\pipeline/store_data_WB [24]), .ip2(n22344), .op(
        n22323) );
  nand3_1 U24946 ( .ip1(n22324), .ip2(n22323), .ip3(n22322), .op(
        dmem_hwdata[24]) );
  nand2_1 U24947 ( .ip1(n22343), .ip2(\pipeline/store_data_WB [9]), .op(n22327) );
  nand2_1 U24948 ( .ip1(\pipeline/store_data_WB [25]), .ip2(n22344), .op(
        n22325) );
  nand3_1 U24949 ( .ip1(n22327), .ip2(n22326), .ip3(n22325), .op(
        dmem_hwdata[25]) );
  nand2_1 U24950 ( .ip1(n22343), .ip2(\pipeline/store_data_WB [10]), .op(
        n22330) );
  nand2_1 U24951 ( .ip1(\pipeline/store_data_WB [26]), .ip2(n22344), .op(
        n22328) );
  nand3_1 U24952 ( .ip1(n22330), .ip2(n22329), .ip3(n22328), .op(
        dmem_hwdata[26]) );
  nand2_1 U24953 ( .ip1(n22343), .ip2(\pipeline/store_data_WB [11]), .op(
        n22333) );
  nand2_1 U24954 ( .ip1(\pipeline/store_data_WB [27]), .ip2(n22344), .op(
        n22331) );
  nand3_1 U24955 ( .ip1(n22333), .ip2(n22332), .ip3(n22331), .op(
        dmem_hwdata[27]) );
  nand2_1 U24956 ( .ip1(n22343), .ip2(\pipeline/store_data_WB [12]), .op(
        n22336) );
  nand2_1 U24957 ( .ip1(\pipeline/store_data_WB [28]), .ip2(n22344), .op(
        n22334) );
  nand3_1 U24958 ( .ip1(n22336), .ip2(n22335), .ip3(n22334), .op(
        dmem_hwdata[28]) );
  nand2_1 U24959 ( .ip1(n22343), .ip2(\pipeline/store_data_WB [13]), .op(
        n22339) );
  nand2_1 U24960 ( .ip1(\pipeline/store_data_WB [29]), .ip2(n22344), .op(
        n22337) );
  nand3_1 U24961 ( .ip1(n22339), .ip2(n22338), .ip3(n22337), .op(
        dmem_hwdata[29]) );
  nand2_1 U24962 ( .ip1(n22343), .ip2(\pipeline/store_data_WB [14]), .op(
        n22342) );
  nand2_1 U24963 ( .ip1(\pipeline/store_data_WB [30]), .ip2(n22344), .op(
        n22340) );
  nand3_1 U24964 ( .ip1(n22342), .ip2(n22341), .ip3(n22340), .op(
        dmem_hwdata[30]) );
  nand2_1 U24965 ( .ip1(n22343), .ip2(\pipeline/store_data_WB [15]), .op(
        n22347) );
  nand2_1 U24966 ( .ip1(\pipeline/store_data_WB [31]), .ip2(n22344), .op(
        n22345) );
  nand3_1 U24967 ( .ip1(n22347), .ip2(n22346), .ip3(n22345), .op(
        dmem_hwdata[31]) );
  nor2_1 U24968 ( .ip1(htif_pcr_req_valid), .ip2(htif_pcr_resp_valid), .op(
        n22348) );
  not_ab_or_c_or_d U24969 ( .ip1(htif_pcr_resp_valid), .ip2(
        htif_pcr_resp_ready), .ip3(htif_reset), .ip4(n22348), .op(n10139) );
  nand2_1 U24970 ( .ip1(\pipeline/csr/mie [0]), .ip2(n22356), .op(n22350) );
  nand2_1 U24971 ( .ip1(n22357), .ip2(n22377), .op(n22349) );
  nand2_1 U24972 ( .ip1(n22350), .ip2(n22349), .op(n10060) );
  nand2_1 U24973 ( .ip1(\pipeline/csr/mie [2]), .ip2(n22356), .op(n22353) );
  nand2_1 U24974 ( .ip1(n22357), .ip2(n22351), .op(n22352) );
  nand2_1 U24975 ( .ip1(n22353), .ip2(n22352), .op(n10058) );
  nand2_1 U24976 ( .ip1(\pipeline/csr/mie [4]), .ip2(n22356), .op(n22355) );
  nand2_1 U24977 ( .ip1(n22357), .ip2(n22360), .op(n22354) );
  nand2_1 U24978 ( .ip1(n22355), .ip2(n22354), .op(n10056) );
  nand2_1 U24979 ( .ip1(\pipeline/csr/mie [6]), .ip2(n22356), .op(n22359) );
  nand2_1 U24980 ( .ip1(n22357), .ip2(n22364), .op(n22358) );
  nand2_1 U24981 ( .ip1(n22359), .ip2(n22358), .op(n10054) );
  nand2_1 U24982 ( .ip1(\pipeline/csr/mtimecmp [4]), .ip2(n22363), .op(n22362)
         );
  nand2_1 U24983 ( .ip1(n22365), .ip2(n22360), .op(n22361) );
  nand2_1 U24984 ( .ip1(n22362), .ip2(n22361), .op(n10018) );
  nand2_1 U24985 ( .ip1(\pipeline/csr/mtimecmp [6]), .ip2(n22363), .op(n22367)
         );
  nand2_1 U24986 ( .ip1(n22365), .ip2(n22364), .op(n22366) );
  nand2_1 U24987 ( .ip1(n22367), .ip2(n22366), .op(n10016) );
  nor2_1 U24988 ( .ip1(n22368), .ip2(n22371), .op(n22369) );
  not_ab_or_c_or_d U24989 ( .ip1(n22371), .ip2(n22370), .ip3(htif_reset), 
        .ip4(n22369), .op(n10001) );
  nand2_1 U24990 ( .ip1(\pipeline/csr/from_host [0]), .ip2(n22372), .op(n22375) );
  nand2_1 U24991 ( .ip1(n22373), .ip2(n22377), .op(n22374) );
  nand2_1 U24992 ( .ip1(n22375), .ip2(n22374), .op(n9960) );
  nand2_1 U24993 ( .ip1(\pipeline/csr/to_host [0]), .ip2(n22376), .op(n22380)
         );
  nand2_1 U24994 ( .ip1(n22378), .ip2(n22377), .op(n22379) );
  nand2_1 U24995 ( .ip1(n22380), .ip2(n22379), .op(n8772) );
  nand2_1 U24996 ( .ip1(n22476), .ip2(htif_pcr_resp_data[0]), .op(n22385) );
  nand2_1 U24997 ( .ip1(\pipeline/csr/to_host [0]), .ip2(n22477), .op(n22384)
         );
  inv_1 U24998 ( .ip(htif_pcr_req_addr[0]), .op(n22382) );
  nor2_1 U24999 ( .ip1(n22382), .ip2(n22381), .op(n22478) );
  nand2_1 U25000 ( .ip1(\pipeline/csr/from_host [0]), .ip2(n22478), .op(n22383) );
  nand3_1 U25001 ( .ip1(n22385), .ip2(n22384), .ip3(n22383), .op(n8668) );
  nand2_1 U25002 ( .ip1(n22476), .ip2(htif_pcr_resp_data[1]), .op(n22388) );
  nand2_1 U25003 ( .ip1(\pipeline/csr/to_host [1]), .ip2(n22477), .op(n22387)
         );
  nand2_1 U25004 ( .ip1(\pipeline/csr/from_host [1]), .ip2(n22478), .op(n22386) );
  nand3_1 U25005 ( .ip1(n22388), .ip2(n22387), .ip3(n22386), .op(n8667) );
  nand2_1 U25006 ( .ip1(n22476), .ip2(htif_pcr_resp_data[2]), .op(n22391) );
  nand2_1 U25007 ( .ip1(\pipeline/csr/to_host [2]), .ip2(n22477), .op(n22390)
         );
  nand2_1 U25008 ( .ip1(\pipeline/csr/from_host [2]), .ip2(n22478), .op(n22389) );
  nand3_1 U25009 ( .ip1(n22391), .ip2(n22390), .ip3(n22389), .op(n8666) );
  nand2_1 U25010 ( .ip1(n22476), .ip2(htif_pcr_resp_data[3]), .op(n22394) );
  nand2_1 U25011 ( .ip1(\pipeline/csr/to_host [3]), .ip2(n22477), .op(n22393)
         );
  nand2_1 U25012 ( .ip1(\pipeline/csr/from_host [3]), .ip2(n22478), .op(n22392) );
  nand3_1 U25013 ( .ip1(n22394), .ip2(n22393), .ip3(n22392), .op(n8665) );
  nand2_1 U25014 ( .ip1(n22476), .ip2(htif_pcr_resp_data[4]), .op(n22397) );
  nand2_1 U25015 ( .ip1(\pipeline/csr/to_host [4]), .ip2(n22477), .op(n22396)
         );
  nand2_1 U25016 ( .ip1(\pipeline/csr/from_host [4]), .ip2(n22478), .op(n22395) );
  nand3_1 U25017 ( .ip1(n22397), .ip2(n22396), .ip3(n22395), .op(n8664) );
  nand2_1 U25018 ( .ip1(n22476), .ip2(htif_pcr_resp_data[5]), .op(n22400) );
  nand2_1 U25019 ( .ip1(\pipeline/csr/to_host [5]), .ip2(n22477), .op(n22399)
         );
  nand2_1 U25020 ( .ip1(\pipeline/csr/from_host [5]), .ip2(n22478), .op(n22398) );
  nand3_1 U25021 ( .ip1(n22400), .ip2(n22399), .ip3(n22398), .op(n8663) );
  nand2_1 U25022 ( .ip1(n22476), .ip2(htif_pcr_resp_data[6]), .op(n22403) );
  nand2_1 U25023 ( .ip1(\pipeline/csr/to_host [6]), .ip2(n22477), .op(n22402)
         );
  nand2_1 U25024 ( .ip1(\pipeline/csr/from_host [6]), .ip2(n22478), .op(n22401) );
  nand3_1 U25025 ( .ip1(n22403), .ip2(n22402), .ip3(n22401), .op(n8662) );
  nand2_1 U25026 ( .ip1(n22476), .ip2(htif_pcr_resp_data[7]), .op(n22406) );
  nand2_1 U25027 ( .ip1(\pipeline/csr/to_host [7]), .ip2(n22477), .op(n22405)
         );
  nand2_1 U25028 ( .ip1(\pipeline/csr/from_host [7]), .ip2(n22478), .op(n22404) );
  nand3_1 U25029 ( .ip1(n22406), .ip2(n22405), .ip3(n22404), .op(n8661) );
  nand2_1 U25030 ( .ip1(n22476), .ip2(htif_pcr_resp_data[8]), .op(n22409) );
  nand2_1 U25031 ( .ip1(\pipeline/csr/to_host [8]), .ip2(n22477), .op(n22408)
         );
  nand2_1 U25032 ( .ip1(\pipeline/csr/from_host [8]), .ip2(n22478), .op(n22407) );
  nand3_1 U25033 ( .ip1(n22409), .ip2(n22408), .ip3(n22407), .op(n8660) );
  nand2_1 U25034 ( .ip1(n22476), .ip2(htif_pcr_resp_data[9]), .op(n22412) );
  nand2_1 U25035 ( .ip1(\pipeline/csr/to_host [9]), .ip2(n22477), .op(n22411)
         );
  nand2_1 U25036 ( .ip1(\pipeline/csr/from_host [9]), .ip2(n22478), .op(n22410) );
  nand3_1 U25037 ( .ip1(n22412), .ip2(n22411), .ip3(n22410), .op(n8659) );
  nand2_1 U25038 ( .ip1(n22476), .ip2(htif_pcr_resp_data[10]), .op(n22415) );
  nand2_1 U25039 ( .ip1(\pipeline/csr/to_host [10]), .ip2(n22477), .op(n22414)
         );
  nand2_1 U25040 ( .ip1(\pipeline/csr/from_host [10]), .ip2(n22478), .op(
        n22413) );
  nand3_1 U25041 ( .ip1(n22415), .ip2(n22414), .ip3(n22413), .op(n8658) );
  nand2_1 U25042 ( .ip1(n22476), .ip2(htif_pcr_resp_data[11]), .op(n22418) );
  nand2_1 U25043 ( .ip1(\pipeline/csr/to_host [11]), .ip2(n22477), .op(n22417)
         );
  nand2_1 U25044 ( .ip1(\pipeline/csr/from_host [11]), .ip2(n22478), .op(
        n22416) );
  nand3_1 U25045 ( .ip1(n22418), .ip2(n22417), .ip3(n22416), .op(n8657) );
  nand2_1 U25046 ( .ip1(n22476), .ip2(htif_pcr_resp_data[12]), .op(n22421) );
  nand2_1 U25047 ( .ip1(\pipeline/csr/to_host [12]), .ip2(n22477), .op(n22420)
         );
  nand2_1 U25048 ( .ip1(\pipeline/csr/from_host [12]), .ip2(n22478), .op(
        n22419) );
  nand3_1 U25049 ( .ip1(n22421), .ip2(n22420), .ip3(n22419), .op(n8656) );
  nand2_1 U25050 ( .ip1(n22476), .ip2(htif_pcr_resp_data[13]), .op(n22424) );
  nand2_1 U25051 ( .ip1(\pipeline/csr/to_host [13]), .ip2(n22477), .op(n22423)
         );
  nand2_1 U25052 ( .ip1(\pipeline/csr/from_host [13]), .ip2(n22478), .op(
        n22422) );
  nand3_1 U25053 ( .ip1(n22424), .ip2(n22423), .ip3(n22422), .op(n8655) );
  nand2_1 U25054 ( .ip1(n22476), .ip2(htif_pcr_resp_data[14]), .op(n22427) );
  nand2_1 U25055 ( .ip1(\pipeline/csr/to_host [14]), .ip2(n22477), .op(n22426)
         );
  nand2_1 U25056 ( .ip1(\pipeline/csr/from_host [14]), .ip2(n22478), .op(
        n22425) );
  nand3_1 U25057 ( .ip1(n22427), .ip2(n22426), .ip3(n22425), .op(n8654) );
  nand2_1 U25058 ( .ip1(n22476), .ip2(htif_pcr_resp_data[15]), .op(n22430) );
  nand2_1 U25059 ( .ip1(\pipeline/csr/to_host [15]), .ip2(n22477), .op(n22429)
         );
  nand2_1 U25060 ( .ip1(\pipeline/csr/from_host [15]), .ip2(n22478), .op(
        n22428) );
  nand3_1 U25061 ( .ip1(n22430), .ip2(n22429), .ip3(n22428), .op(n8653) );
  nand2_1 U25062 ( .ip1(n22476), .ip2(htif_pcr_resp_data[16]), .op(n22433) );
  nand2_1 U25063 ( .ip1(\pipeline/csr/to_host [16]), .ip2(n22477), .op(n22432)
         );
  nand2_1 U25064 ( .ip1(\pipeline/csr/from_host [16]), .ip2(n22478), .op(
        n22431) );
  nand3_1 U25065 ( .ip1(n22433), .ip2(n22432), .ip3(n22431), .op(n8652) );
  nand2_1 U25066 ( .ip1(n22476), .ip2(htif_pcr_resp_data[17]), .op(n22436) );
  nand2_1 U25067 ( .ip1(\pipeline/csr/to_host [17]), .ip2(n22477), .op(n22435)
         );
  nand2_1 U25068 ( .ip1(\pipeline/csr/from_host [17]), .ip2(n22478), .op(
        n22434) );
  nand3_1 U25069 ( .ip1(n22436), .ip2(n22435), .ip3(n22434), .op(n8651) );
  nand2_1 U25070 ( .ip1(n22476), .ip2(htif_pcr_resp_data[18]), .op(n22439) );
  nand2_1 U25071 ( .ip1(\pipeline/csr/to_host [18]), .ip2(n22477), .op(n22438)
         );
  nand2_1 U25072 ( .ip1(\pipeline/csr/from_host [18]), .ip2(n22478), .op(
        n22437) );
  nand3_1 U25073 ( .ip1(n22439), .ip2(n22438), .ip3(n22437), .op(n8650) );
  nand2_1 U25074 ( .ip1(n22476), .ip2(htif_pcr_resp_data[19]), .op(n22442) );
  nand2_1 U25075 ( .ip1(\pipeline/csr/to_host [19]), .ip2(n22477), .op(n22441)
         );
  nand2_1 U25076 ( .ip1(\pipeline/csr/from_host [19]), .ip2(n22478), .op(
        n22440) );
  nand3_1 U25077 ( .ip1(n22442), .ip2(n22441), .ip3(n22440), .op(n8649) );
  nand2_1 U25078 ( .ip1(n22476), .ip2(htif_pcr_resp_data[20]), .op(n22445) );
  nand2_1 U25079 ( .ip1(\pipeline/csr/to_host [20]), .ip2(n22477), .op(n22444)
         );
  nand2_1 U25080 ( .ip1(\pipeline/csr/from_host [20]), .ip2(n22478), .op(
        n22443) );
  nand3_1 U25081 ( .ip1(n22445), .ip2(n22444), .ip3(n22443), .op(n8648) );
  nand2_1 U25082 ( .ip1(n22476), .ip2(htif_pcr_resp_data[21]), .op(n22448) );
  nand2_1 U25083 ( .ip1(\pipeline/csr/to_host [21]), .ip2(n22477), .op(n22447)
         );
  nand2_1 U25084 ( .ip1(\pipeline/csr/from_host [21]), .ip2(n22478), .op(
        n22446) );
  nand3_1 U25085 ( .ip1(n22448), .ip2(n22447), .ip3(n22446), .op(n8647) );
  nand2_1 U25086 ( .ip1(n22476), .ip2(htif_pcr_resp_data[22]), .op(n22451) );
  nand2_1 U25087 ( .ip1(\pipeline/csr/to_host [22]), .ip2(n22477), .op(n22450)
         );
  nand2_1 U25088 ( .ip1(\pipeline/csr/from_host [22]), .ip2(n22478), .op(
        n22449) );
  nand3_1 U25089 ( .ip1(n22451), .ip2(n22450), .ip3(n22449), .op(n8646) );
  nand2_1 U25090 ( .ip1(n22476), .ip2(htif_pcr_resp_data[23]), .op(n22454) );
  nand2_1 U25091 ( .ip1(\pipeline/csr/to_host [23]), .ip2(n22477), .op(n22453)
         );
  nand2_1 U25092 ( .ip1(\pipeline/csr/from_host [23]), .ip2(n22478), .op(
        n22452) );
  nand3_1 U25093 ( .ip1(n22454), .ip2(n22453), .ip3(n22452), .op(n8645) );
  nand2_1 U25094 ( .ip1(n22476), .ip2(htif_pcr_resp_data[24]), .op(n22457) );
  nand2_1 U25095 ( .ip1(\pipeline/csr/to_host [24]), .ip2(n22477), .op(n22456)
         );
  nand2_1 U25096 ( .ip1(\pipeline/csr/from_host [24]), .ip2(n22478), .op(
        n22455) );
  nand3_1 U25097 ( .ip1(n22457), .ip2(n22456), .ip3(n22455), .op(n8644) );
  nand2_1 U25098 ( .ip1(n22476), .ip2(htif_pcr_resp_data[25]), .op(n22460) );
  nand2_1 U25099 ( .ip1(\pipeline/csr/to_host [25]), .ip2(n22477), .op(n22459)
         );
  nand2_1 U25100 ( .ip1(\pipeline/csr/from_host [25]), .ip2(n22478), .op(
        n22458) );
  nand3_1 U25101 ( .ip1(n22460), .ip2(n22459), .ip3(n22458), .op(n8643) );
  nand2_1 U25102 ( .ip1(n22476), .ip2(htif_pcr_resp_data[26]), .op(n22463) );
  nand2_1 U25103 ( .ip1(\pipeline/csr/to_host [26]), .ip2(n22477), .op(n22462)
         );
  nand2_1 U25104 ( .ip1(\pipeline/csr/from_host [26]), .ip2(n22478), .op(
        n22461) );
  nand3_1 U25105 ( .ip1(n22463), .ip2(n22462), .ip3(n22461), .op(n8642) );
  nand2_1 U25106 ( .ip1(n22476), .ip2(htif_pcr_resp_data[27]), .op(n22466) );
  nand2_1 U25107 ( .ip1(\pipeline/csr/to_host [27]), .ip2(n22477), .op(n22465)
         );
  nand2_1 U25108 ( .ip1(\pipeline/csr/from_host [27]), .ip2(n22478), .op(
        n22464) );
  nand3_1 U25109 ( .ip1(n22466), .ip2(n22465), .ip3(n22464), .op(n8641) );
  nand2_1 U25110 ( .ip1(n22476), .ip2(htif_pcr_resp_data[28]), .op(n22469) );
  nand2_1 U25111 ( .ip1(\pipeline/csr/to_host [28]), .ip2(n22477), .op(n22468)
         );
  nand2_1 U25112 ( .ip1(\pipeline/csr/from_host [28]), .ip2(n22478), .op(
        n22467) );
  nand3_1 U25113 ( .ip1(n22469), .ip2(n22468), .ip3(n22467), .op(n8640) );
  nand2_1 U25114 ( .ip1(n22476), .ip2(htif_pcr_resp_data[29]), .op(n22472) );
  nand2_1 U25115 ( .ip1(\pipeline/csr/to_host [29]), .ip2(n22477), .op(n22471)
         );
  nand2_1 U25116 ( .ip1(\pipeline/csr/from_host [29]), .ip2(n22478), .op(
        n22470) );
  nand3_1 U25117 ( .ip1(n22472), .ip2(n22471), .ip3(n22470), .op(n8639) );
  nand2_1 U25118 ( .ip1(n22476), .ip2(htif_pcr_resp_data[30]), .op(n22475) );
  nand2_1 U25119 ( .ip1(\pipeline/csr/to_host [30]), .ip2(n22477), .op(n22474)
         );
  nand2_1 U25120 ( .ip1(\pipeline/csr/from_host [30]), .ip2(n22478), .op(
        n22473) );
  nand3_1 U25121 ( .ip1(n22475), .ip2(n22474), .ip3(n22473), .op(n8638) );
  nand2_1 U25122 ( .ip1(n22476), .ip2(htif_pcr_resp_data[31]), .op(n22481) );
  nand2_1 U25123 ( .ip1(\pipeline/csr/to_host [31]), .ip2(n22477), .op(n22480)
         );
  nand2_1 U25124 ( .ip1(\pipeline/csr/from_host [31]), .ip2(n22478), .op(
        n22479) );
  nand3_1 U25125 ( .ip1(n22481), .ip2(n22480), .ip3(n22479), .op(n8637) );
  nor2_1 U25126 ( .ip1(\pipeline/md_resp_result [31]), .ip2(n22482), .op(
        n22486) );
  nor2_1 U25127 ( .ip1(n22486), .ip2(n22485), .op(n22483) );
  nor2_1 U25128 ( .ip1(\pipeline/md/b [32]), .ip2(n22483), .op(n22494) );
  nor3_1 U25129 ( .ip1(n22486), .ip2(n22485), .ip3(n22484), .op(n22492) );
  or2_1 U25130 ( .ip1(n22494), .ip2(n22492), .op(n22487) );
  or3_1 U25131 ( .ip1(\pipeline/md/result [32]), .ip2(n22755), .ip3(n22487), 
        .op(n22491) );
  nand2_1 U25132 ( .ip1(n14765), .ip2(n22487), .op(n22488) );
  nand2_1 U25133 ( .ip1(n22738), .ip2(n22488), .op(n22489) );
  nand2_1 U25134 ( .ip1(\pipeline/md/result [32]), .ip2(n22489), .op(n22490)
         );
  nand2_1 U25135 ( .ip1(n22491), .ip2(n22490), .op(n8602) );
  nor2_1 U25136 ( .ip1(\pipeline/md/result [32]), .ip2(n22492), .op(n22493) );
  nor2_1 U25137 ( .ip1(n22494), .ip2(n22493), .op(n22497) );
  inv_1 U25138 ( .ip(n22497), .op(n22496) );
  nor2_1 U25139 ( .ip1(n22496), .ip2(n22495), .op(n22499) );
  nor2_1 U25140 ( .ip1(\pipeline/md/result [33]), .ip2(n22499), .op(n22505) );
  nor2_1 U25141 ( .ip1(\pipeline/md/b [33]), .ip2(n22497), .op(n22506) );
  inv_1 U25142 ( .ip(n22506), .op(n22498) );
  nand3_1 U25143 ( .ip1(n22505), .ip2(n22750), .ip3(n22498), .op(n22504) );
  or2_1 U25144 ( .ip1(n22506), .ip2(n22499), .op(n22500) );
  nand2_1 U25145 ( .ip1(n21440), .ip2(n22500), .op(n22501) );
  nand2_1 U25146 ( .ip1(n22738), .ip2(n22501), .op(n22502) );
  nand2_1 U25147 ( .ip1(\pipeline/md/result [33]), .ip2(n22502), .op(n22503)
         );
  nand2_1 U25148 ( .ip1(n22504), .ip2(n22503), .op(n8601) );
  nor2_1 U25149 ( .ip1(n22506), .ip2(n22505), .op(n22507) );
  nor2_1 U25150 ( .ip1(\pipeline/md/b [34]), .ip2(n22507), .op(n22515) );
  and2_1 U25151 ( .ip1(n22507), .ip2(\pipeline/md/b [34]), .op(n22513) );
  or2_1 U25152 ( .ip1(n22515), .ip2(n22513), .op(n22508) );
  nand2_1 U25153 ( .ip1(n20310), .ip2(n22508), .op(n22509) );
  nand2_1 U25154 ( .ip1(n22738), .ip2(n22509), .op(n22512) );
  nor3_1 U25155 ( .ip1(n22515), .ip2(n22513), .ip3(n22755), .op(n22511) );
  mux2_1 U25156 ( .ip1(n22512), .ip2(n22511), .s(n22510), .op(n8600) );
  nor2_1 U25157 ( .ip1(n22513), .ip2(\pipeline/md/result [34]), .op(n22514) );
  nor2_1 U25158 ( .ip1(n22515), .ip2(n22514), .op(n22516) );
  nor2_1 U25159 ( .ip1(\pipeline/md/b [35]), .ip2(n22516), .op(n22524) );
  and2_1 U25160 ( .ip1(n22516), .ip2(\pipeline/md/b [35]), .op(n22522) );
  or2_1 U25161 ( .ip1(n22524), .ip2(n22522), .op(n22517) );
  nand2_1 U25162 ( .ip1(n14765), .ip2(n22517), .op(n22518) );
  nand2_1 U25163 ( .ip1(n22738), .ip2(n22518), .op(n22521) );
  nor3_1 U25164 ( .ip1(n22524), .ip2(n22522), .ip3(n22755), .op(n22520) );
  mux2_1 U25165 ( .ip1(n22521), .ip2(n22520), .s(n22519), .op(n8599) );
  nor2_1 U25166 ( .ip1(n22522), .ip2(\pipeline/md/result [35]), .op(n22523) );
  nor2_1 U25167 ( .ip1(n22524), .ip2(n22523), .op(n22525) );
  or2_1 U25168 ( .ip1(\pipeline/md/b [36]), .ip2(n22525), .op(n22534) );
  nand2_1 U25169 ( .ip1(\pipeline/md/b [36]), .ip2(n22525), .op(n22527) );
  and2_1 U25170 ( .ip1(n22526), .ip2(n22527), .op(n22533) );
  nand3_1 U25171 ( .ip1(n22534), .ip2(n22750), .ip3(n22533), .op(n22532) );
  nand2_1 U25172 ( .ip1(n22534), .ip2(n22527), .op(n22528) );
  nand2_1 U25173 ( .ip1(n14765), .ip2(n22528), .op(n22529) );
  nand2_1 U25174 ( .ip1(n22738), .ip2(n22529), .op(n22530) );
  nand2_1 U25175 ( .ip1(\pipeline/md/result [36]), .ip2(n22530), .op(n22531)
         );
  nand2_1 U25176 ( .ip1(n22532), .ip2(n22531), .op(n8598) );
  inv_1 U25177 ( .ip(n22533), .op(n22535) );
  nand2_1 U25178 ( .ip1(n22535), .ip2(n22534), .op(n22540) );
  xor2_1 U25179 ( .ip1(\pipeline/md/b [37]), .ip2(n22542), .op(n22536) );
  xor2_1 U25180 ( .ip1(n22540), .ip2(n22536), .op(n22537) );
  nand2_1 U25181 ( .ip1(n22750), .ip2(n22537), .op(n22539) );
  inv_1 U25182 ( .ip(n22738), .op(n22753) );
  nand2_1 U25183 ( .ip1(\pipeline/md/result [37]), .ip2(n22753), .op(n22538)
         );
  nand2_1 U25184 ( .ip1(n22539), .ip2(n22538), .op(n8597) );
  nor2_1 U25185 ( .ip1(\pipeline/md/b [37]), .ip2(\pipeline/md/result [37]), 
        .op(n22541) );
  nor2_1 U25186 ( .ip1(n22541), .ip2(n22540), .op(n22545) );
  nor2_1 U25187 ( .ip1(n22543), .ip2(n22542), .op(n22544) );
  nor2_1 U25188 ( .ip1(n22545), .ip2(n22544), .op(n22551) );
  xor2_1 U25189 ( .ip1(\pipeline/md/b [38]), .ip2(n22552), .op(n22546) );
  xor2_1 U25190 ( .ip1(n22551), .ip2(n22546), .op(n22547) );
  nand2_1 U25191 ( .ip1(n22750), .ip2(n22547), .op(n22549) );
  nand2_1 U25192 ( .ip1(\pipeline/md/result [38]), .ip2(n22753), .op(n22548)
         );
  nand2_1 U25193 ( .ip1(n22549), .ip2(n22548), .op(n8596) );
  nor2_1 U25194 ( .ip1(\pipeline/md/b [38]), .ip2(\pipeline/md/result [38]), 
        .op(n22550) );
  nor2_1 U25195 ( .ip1(n22551), .ip2(n22550), .op(n22555) );
  nor2_1 U25196 ( .ip1(n22553), .ip2(n22552), .op(n22554) );
  nor2_1 U25197 ( .ip1(n22555), .ip2(n22554), .op(n22562) );
  xor2_1 U25198 ( .ip1(\pipeline/md/b [39]), .ip2(n22562), .op(n22557) );
  nand2_1 U25199 ( .ip1(n21440), .ip2(n22557), .op(n22556) );
  nand2_1 U25200 ( .ip1(n22738), .ip2(n22556), .op(n22560) );
  nor2_1 U25201 ( .ip1(n22557), .ip2(n22755), .op(n22559) );
  mux2_1 U25202 ( .ip1(n22560), .ip2(n22559), .s(n22558), .op(n8595) );
  nand2_1 U25203 ( .ip1(\pipeline/md/b [39]), .ip2(\pipeline/md/result [39]), 
        .op(n22564) );
  nor2_1 U25204 ( .ip1(\pipeline/md/b [39]), .ip2(\pipeline/md/result [39]), 
        .op(n22561) );
  or2_1 U25205 ( .ip1(n22562), .ip2(n22561), .op(n22563) );
  nand2_1 U25206 ( .ip1(n22564), .ip2(n22563), .op(n22568) );
  nand2_1 U25207 ( .ip1(n22750), .ip2(n22565), .op(n22567) );
  nand2_1 U25208 ( .ip1(\pipeline/md/result [40]), .ip2(n22753), .op(n22566)
         );
  nand2_1 U25209 ( .ip1(n22567), .ip2(n22566), .op(n8594) );
  fulladder U25210 ( .a(\pipeline/md/b [40]), .b(\pipeline/md/result [40]), 
        .ci(n22568), .co(n22572), .s(n22565) );
  nand2_1 U25211 ( .ip1(n22750), .ip2(n22569), .op(n22571) );
  nand2_1 U25212 ( .ip1(\pipeline/md/result [41]), .ip2(n22753), .op(n22570)
         );
  nand2_1 U25213 ( .ip1(n22571), .ip2(n22570), .op(n8593) );
  fulladder U25214 ( .a(\pipeline/md/b [41]), .b(\pipeline/md/result [41]), 
        .ci(n22572), .co(n22576), .s(n22569) );
  nand2_1 U25215 ( .ip1(n22750), .ip2(n22573), .op(n22575) );
  nand2_1 U25216 ( .ip1(\pipeline/md/result [42]), .ip2(n22753), .op(n22574)
         );
  nand2_1 U25217 ( .ip1(n22575), .ip2(n22574), .op(n8592) );
  fulladder U25218 ( .a(\pipeline/md/b [42]), .b(\pipeline/md/result [42]), 
        .ci(n22576), .co(n22580), .s(n22573) );
  nand2_1 U25219 ( .ip1(n22750), .ip2(n22577), .op(n22579) );
  nand2_1 U25220 ( .ip1(\pipeline/md/result [43]), .ip2(n22753), .op(n22578)
         );
  nand2_1 U25221 ( .ip1(n22579), .ip2(n22578), .op(n8591) );
  fulladder U25222 ( .a(\pipeline/md/b [43]), .b(\pipeline/md/result [43]), 
        .ci(n22580), .co(n22581), .s(n22577) );
  or2_1 U25223 ( .ip1(\pipeline/md/b [44]), .ip2(n22581), .op(n22590) );
  nand2_1 U25224 ( .ip1(\pipeline/md/b [44]), .ip2(n22581), .op(n22587) );
  nand2_1 U25225 ( .ip1(n22590), .ip2(n22587), .op(n22582) );
  nand2_1 U25226 ( .ip1(n20310), .ip2(n22582), .op(n22583) );
  nand2_1 U25227 ( .ip1(n22738), .ip2(n22583), .op(n22584) );
  nand2_1 U25228 ( .ip1(n22584), .ip2(\pipeline/md/result [44]), .op(n22586)
         );
  nand4_1 U25229 ( .ip1(n22750), .ip2(n22590), .ip3(n22588), .ip4(n22587), 
        .op(n22585) );
  nand2_1 U25230 ( .ip1(n22586), .ip2(n22585), .op(n8590) );
  inv_1 U25231 ( .ip(\pipeline/md/result [45]), .op(n22589) );
  nand2_1 U25232 ( .ip1(n22588), .ip2(n22587), .op(n22591) );
  nand3_1 U25233 ( .ip1(\pipeline/md/b [45]), .ip2(n22591), .ip3(n22590), .op(
        n22594) );
  nand2_1 U25234 ( .ip1(n22589), .ip2(n22594), .op(n22600) );
  inv_1 U25235 ( .ip(n22600), .op(n22603) );
  inv_1 U25236 ( .ip(\pipeline/md/b [45]), .op(n22593) );
  nand2_1 U25237 ( .ip1(n22591), .ip2(n22590), .op(n22592) );
  nand2_1 U25238 ( .ip1(n22593), .ip2(n22592), .op(n22601) );
  nand3_1 U25239 ( .ip1(n22603), .ip2(n22750), .ip3(n22601), .op(n22599) );
  nand2_1 U25240 ( .ip1(n22594), .ip2(n22601), .op(n22595) );
  nand2_1 U25241 ( .ip1(n22595), .ip2(n22750), .op(n22596) );
  nand2_1 U25242 ( .ip1(n22596), .ip2(n22738), .op(n22597) );
  nand2_1 U25243 ( .ip1(\pipeline/md/result [45]), .ip2(n22597), .op(n22598)
         );
  nand2_1 U25244 ( .ip1(n22599), .ip2(n22598), .op(n8589) );
  nand3_1 U25245 ( .ip1(\pipeline/md/b [46]), .ip2(n22600), .ip3(n22601), .op(
        n22613) );
  inv_1 U25246 ( .ip(n22601), .op(n22602) );
  nor2_1 U25247 ( .ip1(n22603), .ip2(n22602), .op(n22604) );
  nor2_1 U25248 ( .ip1(\pipeline/md/b [46]), .ip2(n22604), .op(n22610) );
  inv_1 U25249 ( .ip(n22610), .op(n22605) );
  nand2_1 U25250 ( .ip1(n22613), .ip2(n22605), .op(n22607) );
  nand2_1 U25251 ( .ip1(n21440), .ip2(n22607), .op(n22606) );
  nand2_1 U25252 ( .ip1(n22738), .ip2(n22606), .op(n22609) );
  nor2_1 U25253 ( .ip1(n22755), .ip2(n22607), .op(n22608) );
  mux2_1 U25254 ( .ip1(n22609), .ip2(n22608), .s(n22611), .op(n8588) );
  nor2_1 U25255 ( .ip1(n22738), .ip2(n22618), .op(n22617) );
  or2_1 U25256 ( .ip1(n22611), .ip2(n22610), .op(n22612) );
  nand2_1 U25257 ( .ip1(n22613), .ip2(n22612), .op(n22621) );
  xor2_1 U25258 ( .ip1(\pipeline/md/b [47]), .ip2(n22618), .op(n22614) );
  xor2_1 U25259 ( .ip1(n22621), .ip2(n22614), .op(n22615) );
  nor2_1 U25260 ( .ip1(n22615), .ip2(n22755), .op(n22616) );
  or2_1 U25261 ( .ip1(n22617), .ip2(n22616), .op(n8587) );
  nand2_1 U25262 ( .ip1(n22619), .ip2(n22618), .op(n22620) );
  nand2_1 U25263 ( .ip1(n22621), .ip2(n22620), .op(n22623) );
  nand2_1 U25264 ( .ip1(\pipeline/md/b [47]), .ip2(\pipeline/md/result [47]), 
        .op(n22622) );
  nand2_1 U25265 ( .ip1(n22623), .ip2(n22622), .op(n22631) );
  xor2_1 U25266 ( .ip1(n22629), .ip2(n22631), .op(n22624) );
  nor2_1 U25267 ( .ip1(n22624), .ip2(n22755), .op(n22627) );
  nand2_1 U25268 ( .ip1(n21440), .ip2(n22624), .op(n22625) );
  nand2_1 U25269 ( .ip1(n22738), .ip2(n22625), .op(n22626) );
  mux2_1 U25270 ( .ip1(n22627), .ip2(n22626), .s(\pipeline/md/result [48]), 
        .op(n8586) );
  xor2_1 U25271 ( .ip1(\pipeline/md/b [49]), .ip2(\pipeline/md/result [49]), 
        .op(n22634) );
  inv_1 U25272 ( .ip(\pipeline/md/result [48]), .op(n22628) );
  nand2_1 U25273 ( .ip1(n22629), .ip2(n22628), .op(n22630) );
  nand2_1 U25274 ( .ip1(n22631), .ip2(n22630), .op(n22633) );
  nand2_1 U25275 ( .ip1(\pipeline/md/b [48]), .ip2(\pipeline/md/result [48]), 
        .op(n22632) );
  nand2_1 U25276 ( .ip1(n22633), .ip2(n22632), .op(n22641) );
  xor2_1 U25277 ( .ip1(n22634), .ip2(n22641), .op(n22635) );
  nand2_1 U25278 ( .ip1(n22750), .ip2(n22635), .op(n22637) );
  nand2_1 U25279 ( .ip1(\pipeline/md/result [49]), .ip2(n22753), .op(n22636)
         );
  nand2_1 U25280 ( .ip1(n22637), .ip2(n22636), .op(n8585) );
  inv_1 U25281 ( .ip(\pipeline/md/b [49]), .op(n22639) );
  nand2_1 U25282 ( .ip1(n22639), .ip2(n22638), .op(n22640) );
  nand2_1 U25283 ( .ip1(n22641), .ip2(n22640), .op(n22643) );
  nand2_1 U25284 ( .ip1(\pipeline/md/b [49]), .ip2(\pipeline/md/result [49]), 
        .op(n22642) );
  nand2_1 U25285 ( .ip1(n22643), .ip2(n22642), .op(n22649) );
  xor2_1 U25286 ( .ip1(n22650), .ip2(n22649), .op(n22644) );
  nor2_1 U25287 ( .ip1(n22644), .ip2(n22755), .op(n22647) );
  nand2_1 U25288 ( .ip1(n20310), .ip2(n22644), .op(n22645) );
  nand2_1 U25289 ( .ip1(n22738), .ip2(n22645), .op(n22646) );
  mux2_1 U25290 ( .ip1(n22647), .ip2(n22646), .s(\pipeline/md/result [50]), 
        .op(n8584) );
  xor2_1 U25291 ( .ip1(\pipeline/md/b [51]), .ip2(\pipeline/md/result [51]), 
        .op(n22654) );
  nand2_1 U25292 ( .ip1(n22651), .ip2(n22650), .op(n22648) );
  nand2_1 U25293 ( .ip1(n22649), .ip2(n22648), .op(n22653) );
  or2_1 U25294 ( .ip1(n22651), .ip2(n22650), .op(n22652) );
  nand2_1 U25295 ( .ip1(n22653), .ip2(n22652), .op(n22659) );
  xor2_1 U25296 ( .ip1(n22654), .ip2(n22659), .op(n22655) );
  nand2_1 U25297 ( .ip1(n22750), .ip2(n22655), .op(n22657) );
  nand2_1 U25298 ( .ip1(\pipeline/md/result [51]), .ip2(n22753), .op(n22656)
         );
  nand2_1 U25299 ( .ip1(n22657), .ip2(n22656), .op(n8583) );
  or2_1 U25300 ( .ip1(\pipeline/md/b [51]), .ip2(\pipeline/md/result [51]), 
        .op(n22658) );
  nand2_1 U25301 ( .ip1(n22659), .ip2(n22658), .op(n22661) );
  nand2_1 U25302 ( .ip1(\pipeline/md/b [51]), .ip2(\pipeline/md/result [51]), 
        .op(n22660) );
  nand2_1 U25303 ( .ip1(n22661), .ip2(n22660), .op(n22662) );
  nor2_1 U25304 ( .ip1(\pipeline/md/b [52]), .ip2(n22662), .op(n22674) );
  nand2_1 U25305 ( .ip1(\pipeline/md/b [52]), .ip2(n22662), .op(n22663) );
  nand2_1 U25306 ( .ip1(n22669), .ip2(n22663), .op(n22672) );
  nor3_1 U25307 ( .ip1(n22674), .ip2(n22672), .ip3(n22755), .op(n22671) );
  inv_1 U25308 ( .ip(n22663), .op(n22664) );
  nor2_1 U25309 ( .ip1(n22674), .ip2(n22664), .op(n22666) );
  nor2_1 U25310 ( .ip1(n22666), .ip2(n22665), .op(n22667) );
  nor2_1 U25311 ( .ip1(n22667), .ip2(n22753), .op(n22668) );
  nor2_1 U25312 ( .ip1(n22669), .ip2(n22668), .op(n22670) );
  or2_1 U25313 ( .ip1(n22671), .ip2(n22670), .op(n8582) );
  inv_1 U25314 ( .ip(n22672), .op(n22673) );
  nor2_1 U25315 ( .ip1(n22674), .ip2(n22673), .op(n22682) );
  xor2_1 U25316 ( .ip1(\pipeline/md/b [53]), .ip2(\pipeline/md/result [53]), 
        .op(n22675) );
  xor2_1 U25317 ( .ip1(n22682), .ip2(n22675), .op(n22676) );
  nand2_1 U25318 ( .ip1(n22750), .ip2(n22676), .op(n22678) );
  nand2_1 U25319 ( .ip1(\pipeline/md/result [53]), .ip2(n22753), .op(n22677)
         );
  nand2_1 U25320 ( .ip1(n22678), .ip2(n22677), .op(n8581) );
  xor2_1 U25321 ( .ip1(\pipeline/md/b [54]), .ip2(\pipeline/md/result [54]), 
        .op(n22685) );
  nand2_1 U25322 ( .ip1(n22680), .ip2(n22679), .op(n22681) );
  nand2_1 U25323 ( .ip1(n22682), .ip2(n22681), .op(n22684) );
  nand2_1 U25324 ( .ip1(\pipeline/md/b [53]), .ip2(\pipeline/md/result [53]), 
        .op(n22683) );
  nand2_1 U25325 ( .ip1(n22684), .ip2(n22683), .op(n22692) );
  xor2_1 U25326 ( .ip1(n22685), .ip2(n22692), .op(n22686) );
  nand2_1 U25327 ( .ip1(n22750), .ip2(n22686), .op(n22688) );
  nand2_1 U25328 ( .ip1(\pipeline/md/result [54]), .ip2(n22753), .op(n22687)
         );
  nand2_1 U25329 ( .ip1(n22688), .ip2(n22687), .op(n8580) );
  inv_1 U25330 ( .ip(\pipeline/md/result [54]), .op(n22689) );
  nand2_1 U25331 ( .ip1(n22690), .ip2(n22689), .op(n22691) );
  nand2_1 U25332 ( .ip1(n22692), .ip2(n22691), .op(n22694) );
  nand2_1 U25333 ( .ip1(\pipeline/md/b [54]), .ip2(\pipeline/md/result [54]), 
        .op(n22693) );
  nand2_1 U25334 ( .ip1(n22694), .ip2(n22693), .op(n22702) );
  xor2_1 U25335 ( .ip1(n22699), .ip2(n22702), .op(n22696) );
  nand2_1 U25336 ( .ip1(n14765), .ip2(n22696), .op(n22695) );
  nand2_1 U25337 ( .ip1(n22738), .ip2(n22695), .op(n22698) );
  nor2_1 U25338 ( .ip1(n22696), .ip2(n22755), .op(n22697) );
  mux2_1 U25339 ( .ip1(n22698), .ip2(n22697), .s(n22700), .op(n8579) );
  nand2_1 U25340 ( .ip1(\pipeline/md/b [55]), .ip2(\pipeline/md/result [55]), 
        .op(n22704) );
  nand2_1 U25341 ( .ip1(n22700), .ip2(n22699), .op(n22701) );
  nand2_1 U25342 ( .ip1(n22702), .ip2(n22701), .op(n22703) );
  nand2_1 U25343 ( .ip1(n22704), .ip2(n22703), .op(n22708) );
  nand2_1 U25344 ( .ip1(n22750), .ip2(n22705), .op(n22707) );
  nand2_1 U25345 ( .ip1(\pipeline/md/result [56]), .ip2(n22753), .op(n22706)
         );
  nand2_1 U25346 ( .ip1(n22707), .ip2(n22706), .op(n8578) );
  fulladder U25347 ( .a(\pipeline/md/b [56]), .b(\pipeline/md/result [56]), 
        .ci(n22708), .co(n22712), .s(n22705) );
  nand2_1 U25348 ( .ip1(n22750), .ip2(n22709), .op(n22711) );
  nand2_1 U25349 ( .ip1(\pipeline/md/result [57]), .ip2(n22753), .op(n22710)
         );
  nand2_1 U25350 ( .ip1(n22711), .ip2(n22710), .op(n8577) );
  fulladder U25351 ( .a(\pipeline/md/b [57]), .b(\pipeline/md/result [57]), 
        .ci(n22712), .co(n22716), .s(n22709) );
  nand2_1 U25352 ( .ip1(n22750), .ip2(n22713), .op(n22715) );
  nand2_1 U25353 ( .ip1(\pipeline/md/result [58]), .ip2(n22753), .op(n22714)
         );
  nand2_1 U25354 ( .ip1(n22715), .ip2(n22714), .op(n8576) );
  nor2_1 U25355 ( .ip1(n22738), .ip2(n22722), .op(n22720) );
  fulladder U25356 ( .a(\pipeline/md/b [58]), .b(\pipeline/md/result [58]), 
        .ci(n22716), .co(n22724), .s(n22713) );
  xor2_1 U25357 ( .ip1(n22724), .ip2(n22722), .op(n22717) );
  xor2_1 U25358 ( .ip1(\pipeline/md/b [59]), .ip2(n22717), .op(n22718) );
  nor2_1 U25359 ( .ip1(n22718), .ip2(n22755), .op(n22719) );
  or2_1 U25360 ( .ip1(n22720), .ip2(n22719), .op(n8575) );
  inv_1 U25361 ( .ip(n22724), .op(n22721) );
  nor2_1 U25362 ( .ip1(n22722), .ip2(n22721), .op(n22723) );
  nor2_1 U25363 ( .ip1(\pipeline/md/b [59]), .ip2(n22723), .op(n22726) );
  nor2_1 U25364 ( .ip1(\pipeline/md/result [59]), .ip2(n22724), .op(n22725) );
  nor2_1 U25365 ( .ip1(n22726), .ip2(n22725), .op(n22732) );
  xor2_1 U25366 ( .ip1(n22732), .ip2(n22734), .op(n22728) );
  nand2_1 U25367 ( .ip1(n14765), .ip2(n22728), .op(n22727) );
  nand2_1 U25368 ( .ip1(n22738), .ip2(n22727), .op(n22730) );
  nor2_1 U25369 ( .ip1(n22755), .ip2(n22728), .op(n22729) );
  mux2_1 U25370 ( .ip1(n22730), .ip2(n22729), .s(n22733), .op(n8574) );
  nor2_1 U25371 ( .ip1(n22734), .ip2(n22733), .op(n22731) );
  or2_1 U25372 ( .ip1(n22732), .ip2(n22731), .op(n22736) );
  nand2_1 U25373 ( .ip1(n22734), .ip2(n22733), .op(n22735) );
  nand2_1 U25374 ( .ip1(n22736), .ip2(n22735), .op(n22742) );
  xor2_1 U25375 ( .ip1(\pipeline/md/b [61]), .ip2(n22742), .op(n22739) );
  nand2_1 U25376 ( .ip1(n21440), .ip2(n22739), .op(n22737) );
  nand2_1 U25377 ( .ip1(n22738), .ip2(n22737), .op(n22741) );
  nor2_1 U25378 ( .ip1(n22755), .ip2(n22739), .op(n22740) );
  mux2_1 U25379 ( .ip1(n22741), .ip2(n22740), .s(n22743), .op(n8573) );
  nor2_1 U25380 ( .ip1(n22742), .ip2(n22744), .op(n22748) );
  or2_1 U25381 ( .ip1(n22742), .ip2(n22743), .op(n22746) );
  or2_1 U25382 ( .ip1(n22744), .ip2(n22743), .op(n22745) );
  nand2_1 U25383 ( .ip1(n22746), .ip2(n22745), .op(n22747) );
  or2_1 U25384 ( .ip1(n22748), .ip2(n22747), .op(n22754) );
  nand2_1 U25385 ( .ip1(n22750), .ip2(n22749), .op(n22752) );
  nand2_1 U25386 ( .ip1(\pipeline/md/result [62]), .ip2(n22753), .op(n22751)
         );
  nand2_1 U25387 ( .ip1(n22752), .ip2(n22751), .op(n8572) );
  and2_1 U25388 ( .ip1(n22753), .ip2(\pipeline/md/result [63]), .op(n22759) );
  fulladder U25389 ( .a(\pipeline/md/result [62]), .b(\pipeline/md/b [62]), 
        .ci(n22754), .co(n22757), .s(n22749) );
  nor2_1 U25390 ( .ip1(\pipeline/md/result [63]), .ip2(n22757), .op(n22756) );
  not_ab_or_c_or_d U25391 ( .ip1(\pipeline/md/result [63]), .ip2(n22757), 
        .ip3(n22756), .ip4(n22755), .op(n22758) );
  or2_1 U25392 ( .ip1(n22759), .ip2(n22758), .op(n8571) );
endmodule

